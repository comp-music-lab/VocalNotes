BZh91AY&SY��%�[6_�py���������� � ��              ��       *��   �           �  7�  Jw��{�����/ܦ� nc���h<$ c�'��6�v�+�%4w�ݎ��xe d-iX���@�y¼Ż�3]ha��5��[�s��)���
PPwt����z�4���G�Pw���L��oC�B�  =�=�ӯvy4ѭ�Xt�!Aq.�OP��u����4ɶ��o^�Ѧ�dx  :X ��xӓ�&��9�:n�d2�pܹ^�r8  7#/N�9qӐ%�-��瓓M4kC¨o  �g��B��hP�C��
(�С��B���(PS�(H  B�*��P � 5O�&U�# F  @i���E?%*J�F�2bi�44��#?L�T��҃@       M��5J���hb �CM &�M$ U(��2�� �ML&�M��I���2=5=&���.����ٍ�"�|�
"��"�DE9)���R���c�������X�I �* �F�{-�U)Om� 71(��* �e*.���\��޼� E?2�����k�x���葹�����ᕳ-�<�)}�Vv&/��I�gH��J�X��ʶ-C��=ѷ7H�xb�t"�����|~�O�����?ȭ��;���g@�<�X,Ґ�������i8N\to>Z7�soI�u'�7u1���E�xį��#p�Sv�_�W�m8&���/�R���w:(@fs��lzJَ�Q��үG;:� ��@���<��p��!	��΢Jݥ�hå�#)b��]�p��P�ܷC�@l^�{'`�]s��z���2/����.{n6t揇�N�cZ�+j�*x2��u��m�>K��7:�ľ�n���lS���ou٥d���g�va��A4=�t�a��ъ������DtUb�cúƍy�M��R�K��EK�<ބW�sO4댜{r�ԧF��1*aBѭ)t���Ö=Aj���pΗ�٤-gC�g.��5	X��������N�K���ء�Lq
T=Jg�T��^r��얎D7On��;{ib�7����������⻏�!ݧ�spҳwm����;�q!��I괍����<s�mg4�tJ+Z2�r���m�pSح܌owX�;C;��k�^���9������^�
u=W\ǳD�m�'X�^�,�
؎�+d0W�=�ծ�����n��cE*�agk�V]���(��cﷸ�9���x��&����zX)�\H�"<���R�E��gcs:.9)�ѯY�b�X��ĐN��z����-�Ɂ$JS�1���8�y�����ś�K<�uT,WDׅ�˸b=��͹V[Nۻ5�����V8��w��� ����S�fhU�ȍ˽�r9j��\1ѧy��-�K{�\�b]Y���>7��y�����+G;s��u�yQB�����3Dy�� ��k��6�±�䖹�9Sܜ�q��3N�s��Y����^@tl�7��K������Z�S��X�n) /a��{^8XS[��Fm���j����e�&�E�#����`�n�xu�M���O/���Z������q����p����`��s���H�9��OA3�G�[ױ����̧˩
[�4��1Q��O0��IH��Y²+��<�BV�]j][�q0C3@�#��!Rx�
}(gk:*���k_l9��&攉$2��u:kw�pSv:c:B�@��cE��8�t`Pnj�{`��$��O��ܝ��%�3�ۖ�S�˻t`�×�f���H�י�d��:��Úb�2ú�����:�=D+�1����	T�Ϸ�I ��ؠ�Bb�Z���vЮV�2~ ���[}.\��4IG�ӰD#�7�G�7�=Ɔ�����*��7_9�k�f%�T8�^I�z_	uZ�<9��0��No�gsq�n�Mu�*�������(� ��곦� [m�w&�Ø�[�A�a\NEf�	��	�頸{�w���QS!�N�v�c5��q�;��L�·
]˻�_b�����8�y˹�!�U٦��xu�B2u�nMػ�v�=��0�� �JR-9��s��>T�2���x��f�roæ:���X����ו��4x��J��՗)��O8��q�Hq�ϯs��Z�pX.P�n��q����7Б�7g1I=-���N��.�@]=���w2����/�)�6v�8�'_kXj'�a8@d}	<�J�?U&��yjܒ^������#s�O�4�z�����&�y	[�^�kPL�IP��SA���-n�'l˹�H��a�p���n��;!uײ'�W��uR�����T>��r#���&XX��'6��#�Gӊ��sk�fh�Qz�7'D��o �r����W!;^�X���g���>#��q�y���7'RwF� ߺ<�69���i}�5�ZW�X$"Ǣm����ƪ퓷�N�r����ze�׫��=O[��w�%&�w�V9ٴE6��g\t��w��L��c�wq�0���kTW��;z�i[w:buRɿ�;�Q�f�r���a�����xFߦ�!�OL�N��ǿ&��ځ��}ܝ��k���v��WP;���*���o.�'b ӁMA9v���ĸVp�hw��M��/X�p�g,|���	�q��n=�sA�N�ثͺ��$,t��-p�efef�d�t��ڲs�r���p�/����+�K�9����R�����v�s��ؒMp�4\�]��j�QZ�=�C�v�ѯ�̼��|7wF�q�н9E�]�s ����W2�4EUr���<��aݙ�N�	P�"��m����d�����L�6hǹݜsbO���@*ƚ�GiL�-ӷz�٬�2s�N5wY�KD�R[w�S��0q��3Oc��g0������"ӌ�/M���5�G����cS�����O5���[u�ouw�4(��<d�M'�Bn�C���:;�"�ٵ(�����N�+{.c&b8�	a!�[#%�J4Y�:|3��噖K�\|[��ߘ�&���k����=�Eus'���!�:8p9�ۗ���£�z[n�(_�_�y��'u���qёU0`�jt�vڪ�.�a��f}���]v`8�닪y�ƹ�Mk���S9;q$���,�u����K���8�iԾj�6A�mS�	4�"�Gma��#6g�<�7;�X;��m�,r/F�7&��,�]e�4M��������Zf��_���iG��SӮӫ�ma ]�mk��;rt�K/�G��]�Ҟ�Ѻzv�á��\�.�mg�R3�&���mk��5ۭs��km��k�s���fո�^�=���B��sv�s�7�����v��A�̕����F�/>-Í�Z�q�v��d5�=''��x�����q���lH�[�t�[f�.�C�����8-6�g�:l6�zl]3Wh��oR�m3��-�dìq[���;�^���n.�;T웓�?]����;�;����0n{7;�֗��wmݽG���ٹ�۵���:.v��vN�[��y݉wX��չ��xqؖ���F���d��s�C8�l����U<y����ENnuW\r�g�;P���F7��s����ͫZF���e�~E׃�
��$8";�(܋�31�9�;fW;u�	�v�m8+#����6+TKśu�Q����O�����
7(�콎؛Yl>�[O]D^z�v[�=��wSim��/[mO�����9�^s�yt���]����\���[V�����������:�玉7��7
�z������G9��i��GN�t�^��t�Ӄ;�׶y���5�wD�g�2����%���F��<y�]���r��\g�������d>�Zܷ�v�̉x��R�c=��'n�W+��u����oZꪮ˜Di���׏c��ɧ�t{e���7o[lp'X��'c:�`h\�y�lxX�k{5��y{�=�٨A�v��;u��W.�J���2&�1��c�z�<���u��<��6�%��JvN��G�/���Ǖ5pg�Y��\��<�v�]�����:��GA��X�wb���k��5úŪ�o]�Gj��}���l��A��U�(�랮��u`k�p�n���A 吠�TdM�k�Qe���xi��2��)z�`��ɩ��ˣ"�mu�wX�۷<V/ͣ�=��g�Ӱ!�m����SO<~>���vk�ݳ[/ ��s6zNƶݍuO.�Z6�py���(M��;W	�.n�:�JS�Rn�I�\n��}�Yx���cv��{a��z���xZ2?�t-C@6�J���9ـy]ml񱞓<��ֱ���-�l�gm�8(q�=qs����z���Z��`�f���Dm��r��ӻ>�;p5�c(�U���+~>��K��j��箭�F�2{b�ɮ5v��Z8���q�1�GeN�q�I��[Wm�ccE�מں)q����p��汛T��M��Tݛ�n�۷��m�����\���h���\��`�<qUŹsP{Y�
����ۧ1v����@�7�덱��*���"b6�-���ם�.���2{'+;{izQ���5������>;�y��t���V�v��n1ss��*a�p絩�X�`�ɥ&����r��3�p�{]�Ϸ+����9y��F��=��mŶ�[�7n���P�����j��W!G0v�g�c���=pi㫎���+��8z��F+���x{8׏Ї�7��AE������aΝ1�gK/�v/<���n|��ltf듟Vk�O`�S�ٸ�P�^<��\vv�v�6�f���g��|F���e�v��.;]�N�vs� ��ՏMOk���ۏ(k�;e�%�����]��mg�ώ\y��5s�w@ܾ�7��m:{;�tl9Ϊ�F�vU��y��m.&�н�(�v�B���ڊ��SeR6]��WY��[�ǣ��� A�u@��I�2�`D:�ľRP[�{y�;�|e��_�+=:su4έ�׉<_��}�����;���I���h���C���1톃w�~H/e�|�TZ��<�9lH�ag������{��bޯ��=;x?�˜���6����,�kD۲�/���ឈ�f�Ƕo#�'j@�����=* �}�$�
x�TV��"�p^�u���ʋ�I�հ,��ôy챸-��=�}�7�b����p�ן޽���l�<�B��τ=)�x��.��R<1cCmk�����;^iTܳ,��=Ӿ��v���}���bh=�åf��x�o`��"kw�&Sۣ�n:���G,�
֗;���Gi$"��Ҳ� M9��o|�
���w@�m6�OI�o�Ϡ�҆��z��{f��#�g^���3���OP����{ٰ��`�;��৹�����
(I����.�Cޱ����F{��a�GM}��7ç7G�������w��n���%���ｰ���vW6��/�)N1�Y����~�{�����erS{ny����ݞ�!��-u��ױ�|0�
]f�{����t�Sj�ˇ�+nh����(��{Ho���/=�ong`^0x�+>q�i�[_��}��H9ވ�>wz3ڄ>�|�K��N��p��{ib}:\�j��a�ƍw����f�蟴,�8���~�@�լ���/�	�Yu��u�uv눟&�3מ��k�u?-��5^[{� �{�Y<=�=�~x���N�zqi��sxd�f��<���W��A�������Ί���x�~��^�.Q�7s��ot�Д�r��G嶺\g��l���hKs�U3n����ێ9��}�F�;>N)�~�!7�1��Ӹ�B2.h���e�����f8��T��"Ѱ1*�lgv�>�q��r�xkCz!�	��ji�^�5������v
���B�y�����p�1omK�������㧰%�O��;];oi��ӓ�N���W1�IW�<�V��jծ>V���:uz8�?�'�o�~ٽ�s=٨﹕�W���_e���.��O�/EN��1�Og�u���<�w;٣NW�\^�5b>|3�C�p[���L�ܧ	�$�;��x��q��MU��5�A��˘�v\7�I��Y�Wv�Jf����G�3���-�����7��4��-Ǜs���.�X�����R�2��P��L=�q�����=���4c
a+��ݎ_.~�>3�4�)�Gt�O������os8�p�{��M��g,��ޜBNO1<�s�x��ڦ�V�tte��݊���ڛd�X������r�;�#I����4ߧ=��O�V����{{ݽ@:�2�z�^�g����'��b�y��l�?G���6���c��V�	s�4[�/��Ƹk0����zϷS�o��dX�5oR�S����nn����Er)�W�E�=�ׇz<j��:!�{"9ޔ�����}�E��p�������;'�y��.�+������E �I���D�.����.m��o�a7n�<}%���<��O۾�_�v88�](����4�����}�({��X���^=�}��k�1��U>?S�;���`}�қ4���Rݙ�;�{녭}�g�<{h���0v�������拓h�\�nn�ىLQs�_v�7k��� �N`���J���ۢ���-��X��q�+�^2c��v�Un>5��ݛ�/{{Nz^�.�Ӽ���I�7���Q�.Jg�I�6/�E��m <���8�o��H�=Fr�n��d��e��"gy{��e�L��y�1fy����P��t?Ts٪:�IA}��eޛ��C	�`�ދ|�s.��+��U����;7֜�1��wg�ך��o�`뻏�i�{��2����ڲ{|����d��k��-�;��cgT�<����n	����ǴU�]��V*��vV����_i,��Nz?n�@S8	�ݏ���-�W|�f�d��<R]û�Ͻ65ZXןdݣ��.]�>���f}��R:�獯!�Ozq����s���i{ϡK�'y�)�s����[XA�2,Im�a��w��9��r���x��&����2��x�/
�["b����fY��*�#Ŵ���!�ȝ{��Dw����ٻ��˹�v�<�]�(���~r�^�p�n<���T��fl�Ǌ���un9^1��r��d��7w���I��:-�ݼ<��uo��D�a�����P1�Ԫ����8�)�^'s���}5{ѹ����N�ʜ��/f�-�n����۞}6�Q�P�~��͡���B˧c�9*��=���8�<^��]��E�}��g@��O[b]�}n����l�m�
�����>�}7��yoaP���sg��{�;��%�����qZ�;��RD֞�J�6�|�R�W��.h������&�{��ۯ`�ڳķ���:{��x�H3�8q[�ʕ��-��Ǘ>s���W����8���Ѭ�g��{��6�R[�'���j��k���3C���{���%��8��0�r�q��;���g�?��fg�}�),%uy~��+��nel�D"cUc��5u��֚&9S��ͺp����.̞�ewYl�2ɷ��L����r/dN�Z|���ls�	���6�q�i��k�u�e��q�s�>��������w<]�u�����퍫�`Y��;-�t{l/]�Ը��;
�z{��nxW�\�y�!v���6��##Ʈ݃���08�=���
�k�u�v����9$�8�c���\��;-���n�\ԏeMԽp�a�j'��v��<Y{9�}�b7\ٺ㞜��V��=a�=��sY�K^����mct;�ʱ�E��gc6��uan�k�V�nu��,�u��Ǌ��G�v��x�dޤ]�֫��sz�6�Um>��7V�9�6T�Dl�U�q �]�>�e�o�{�w���p)�~����u{�\��K3�p�y��7�V	�Oim�n6!��S���ȶ44O;ǆ�1� ���ۓFW�	����7��#�>X1��a���x=%�F~Y~�g���\���$6�m9�BJ�7����уȃO&���[8���E�6|���fˇ�L߀Y~i9�*
fqQ�|HE- |>J�m�M7!�3��9��k9hs'����p`�}0gB�d��9|�p2��'C�񸹙�ka�%�i�Z��hM�rˋ�h�-y��B�6}<Y���k�'���tq�nO��nf{V�Sj���@p�.]pWm����I0��vS%q-�KUL��.c�K��mx�1'�5��v�}<�j.�W_ ��m&Ԍ!�}�SK���׾u	:g�dh��f�_�M��/
��������6��u�u��^w	Q�� �~��5�Z��XMe����4�7վc�=\}�n~x_յo;˳�U#��{�4���w��0��r��Ӯ�'i���>4F� ��
)�j�*X�B�%x��62I[%%+�[��ͯZ����ͬ��^c7�N�G�#O���3g�xɷ33;s�g�m��;b���ھ��3L{g�v�ve�k[ͱ��<���b�'}s�O6� c�p ~ܪOC��|+�$Y�{��g̳ϱ�Tr����7y�	��F���N��'}c��0�88�/`�Oڪ�uIui6��"!<'�;��k��{�X���wn�ُ[��5�kݜ�y�"(�f����9H.z{�G�x�K~�0��r'IDVꩧE.1A[[{���=�~z%~y�0V� �	�~�ƚִ��B���M�Ѳ�
|>;aD��C�4o�2ӊ?a��إ�U����y�5l�~Ӝ���Z�p��p�/��0+V��u
C���댊;az��r����݇�Ȭ���]mμ��[�4P��=[�n�K�n�z^�W�3�����*�b���(:7��.k�Cj��[r8KY[",�%��Qwߐr}�$��l�����/1����6�#L�-Ͼ�>Y�ٓch�my��ړ�f}��<��jCAU �q6�D$Ӏ�<�����7�h�{qlLT�	���ﰛ�� I��7�)��TEAAUT��뫽^�nwn!83f������Kz!'ｯ҆����m&ӑ�_�L��U��䉦�g�:���1����p���5A�,�"�����md�y���0w�Mܡ�����$�6�B���&�.&��ӣ��6�u5�A�Q'�A��B�Vb��V>�U8�4mpR,��W�S�WW�F��a�-1�ˆm������iՙha���s]��V��
�7TO�TF���N�3��t�%��'Z/G��Sp��n�8�9��Y�q��ʈ"�Izצ6��(��TDE"�*,�S�8���o�bZ��B�ә�{�g5h�T+dXX��j�ڌW���d��Ä�w��թ6����Ah0��N����}���Bp\��ׄ�:k�r�z�z!'X��,n�&��=���y�6Ё�D�hY��R��Я�|�@�`X�hx�Y���7��g��s2;�r46��X�wbq����]v�v���fMp�\�hn��F�>x��?[�~�ta�PAb����5vZۻv�lF*Ul��
P���H�O����z���47p|��/4Ѵ2��>���̋�ܧ
��|����@E��[��S�C>��rm�`�^r8��-�@Ad+i���u�|4��>w(h�	����/EyP��.'bf��2�x�y^Vs{Y9A�/(�?�*��V!�<�=�7�0��1�r2�B���>gQ�m����T���d��MF�����|Ey�y�p!��[0XA0ȁ ��e�-֙����C	�m+�W��W>{~�z�3;�O�����^����³F�3�T#�=�3V���6��?�L�w��ߦz34���lҧ{�(�f�ѯ)���޵,2+���zrFlў��:.h�od�Cc������.�a�yp^�llˤf篽���"���[1�^G|@�?���$����,ǲ�Oz�!� ��:}|D�x|�5>{��ʓ�H$���}���5���P�ꋳ���\�uƦ��It!{g��h,����62{|���ˣ�vV{�����O�Z+���q���ZW>��m�ǵ0���7VD��1U*F,��9��!�d݇}���ޞ��q�?��!Dw[�d�N��$��a���0K]�O�_<lh�`�@lV��u�L2L(��O��z.$� �h��*Y���y�^�'JL�k���G;�y�]��%��
O�ߪm遂� �x���>o���0	p(�O�T��y{�.h�^��F��%I21�[���U,������/z篶U�xp����%�4�Pލ�s�O,��Tgò ��C�j�F0	s�Õ\�K⬋K�m߉ѿ7�'G��QF(�o��&0���>�p���ȡ�J�y`c'l*���2�����a\�:3�+��Yr�sLi�B��6,	�lc
�Lj�J�ow�1q��qlK+ŗ}�!5�>�gV>pI+�qI�D4��̖֭�v����ݵ#��������j���tʅ��&�R��l`Z����\�ڃ�� ���y�cUc����"�����޵��~;��Z��OLY��/{��v�Q,d�QH�R�a����W��wd9�I���$������y���Ho�$>��@�y�K~>��L�kE6�ʁ��:"O��)���$t�s<���hw>��2s2AO��1;�a����W˹�C�����4ɿ�1��,�B���|#+��=���ȧ1U��*n��z�QXsO�8�����BmP�*v��[��c{V��vn���n�u�$-�=5ù] t�j3��klK9��;��{gs�,:Ԯ��Oǀ �UUX�b�E���z�����+���a,r�M�x,1&�V'�2�ܐS��^�͡���ܒ�3��M����5���=��껆�2��rN�B�~���Xc|뫟c�w8��}�AO���`�+}�2+kԬ)Q4ڐ��yՆ��f2�2AN�g�{�K�O/a:�coV�Mr*4~=��O�b���_�=���lG�va���A u��]�t}#�}.�w�(�����4����r�lVjUC��k����U`�,AAQ�1`�����<��ěa�2�'��&��~�r���<�B�lg�#��7r�p*}���80��@��;rAOz<>һ�ğwa���<ꆙ�̐Y�$�}=����Әi3k�]<f�~o�C��;��Y^9 ��Y�4��,1?_|��}�="M$�q�c*n2C��t8�AO>�bNn�|����Y��Z���w��髂�J�L�q����H�E��������AE�� e�i}� �÷��s5~JI�SV����A�Y��$v�ֺJ����CT��줎�id+Y���K�.����!�����#�hG��u�w���	���7Ձ�5�="I�z����w.���*J�}}�@�N[ՠw{p���G޽�9��ĝ�a�r�0��$��v�W-d�,�_h�8�/���jS����W��������3�~��J���i����9Ъ��(�(�dA��Eb���Ğr�}�:��:�d��ByNw@7��u8�v�Bm�چT��=���9(��yuc ��o�\"j��u:��]����ulD/�s;l^���ҸʗD �Cm�A�T�}7���\���B}�8AN��c0�9�k�oS�>�o�S�C�0��@�vc!����~Y���s���߽kG��f�k�����2���{�"lW����uԘڗ�qי2�l�M����U��v�oޝ??t^��.ޞ�՛��=-�f�t�7X1К�Gs�us��Lq��֝8EF"E��0QUTAX,QdWC���3Eub�d�ڹ���{��k��p=I�
��vc!��d�aߔ�$v�}��spP>ꇀ 7ے
{Ձ�4Ò2�|�|I���P;�$4��`�y��}��x�.&�vA�/�aI��و���)���𹚁��[� u�4�}~rAO�`bN��<�эp��kIu�慭��];.�݆�>��gV��g�I4��`�k���_3'�?}ˋ�����������p���蚜�!/Vº~�V53��?�$X�*�TYb��UX���g,d��@�vbu"�w�w8.�,��0ݰ^�O�f�_�S�z���n<%$�l1�Y�}i� B��b����to�<�����ί<]�J���+DR"[lV
ǼY��hՅ���=rG�ՑbI�H���'@z�x�(�wRxĚ��������o�9d|�>'y�K��s��zS)���9���f�;��?��QUX,X��,U��H�>�=������tk3~�C���Ts������_"�u\��t ~ŘD�]����P��,cc���*�� �fI�tF��P�,�;�CǾ=>H�c�~�z�������WN�nW�  |�#	xq�W�#��Sg�X�{����|,,�.�3p��ϯ����"	b�!�"�O��޲=:�3&��������<#�vƇY�*e�������T�Hբ�ݓ�_�*�#�N������Ħ,�����Qf��Xx;&�Ӯ.�|��v��������﹏(����xY�i�	��N|���$n�2o;弮 x�d�/j	:�W�2B!���:����
��Νv�o����f�__�4���}k�M�o����ߵ���9%��o	L�äg��	!�&>S�����U�uD,,7Wb�`�2ˆ�_e{��>���bM�P_�l���T�����z�n�+}�#��)�F���8�~=�N�^4�x.�I�7׾>�.N,����:s�笗�.^x�uN���8+پf��_3��#�ד^L/3�<<:�0F�ų�S�xѭ�gn�,�ݺ���W��n�;���W���g3��ssN~_��C���㭸?,7�	���O�ba1�E�ݙ]��z�/3�z�U�l'��!���6��u3��t���U��TQ[4)���"�<E��{$�v�n��u\����"g�V�&��خa�Qmk��C��ډ�1����c�����l\[���l��\�4� �%����v��Xnf�n�=����w�m����
��k��^=0u����9�F��O��'�9zi�x�9\m�]hڸ�y��wZܖ�O�w0�v���+h��]N
�B�B�1�1sV��^�nMq��&��v�3˅���V�լ\}��_?h��{�!��sa��K�8�0#:�Ɨ.�,h�u�8��ܽ��sm'.:zN�g�8؍����v���h1/T�۶�rC�4Y�lVnY6��;�(��z��+ۭ7:'tҙ�bEQ�"E(�"tR��1��.��/Qh@�&V!���	�JP�Χ�����(^h�{�-�dV#��-�c;du0������$�I�" a���{�e� ,�}�Ǧ��]�yޞل�\��Y'B�}���W{x��4� �b?�?u�U�^�����4���E�dv����;�ë߯���l�݊X+}�E�n8y�>�3�tCi�)߯�b3`}�xx$ �P�7l��--L9��x1Y}��x�3\�X�X�k��@�zs����}��o(\�¥�i���l�v9Su��n�߷}��|�^sƩ��)�1�fe�r�sV]]*�AH�
1����
E���y���$Dp��P�j��$�'u�կ}�Gz?Bidm�sퟖo}1'�����G�o2��w��N����F��1%!�>�}��ט,Ļ�}�8�Y���ﾛ��]���2yW�n>R�C�ǝ'j�WSE��5&5+3y�SZ��O�w�3M��}�f>����fO[U�Pz1F�>��⨄j����h�j�[�og�y���γ��,"����
E�DG��){�1�>�@��t|g�8���2�W�f.�w�(,M��� 6ᚴΥ��|>����~`��͕�G�M�n�������9�:;rGI�㻻���,s��j��(I�-}<~�3{~��BJ�-���/ @���<� ����	��?0FG-��"��ĝzehU��_w�w���9�l`��UF,AP�	�w�T�׍���ߠ�/�\}�[�Y���6.�|�{u��y�_|������"�B����b��V�8�-X֖������fa�>	��6�w��U,���Ą�(��x�aV��w����f*�#�y��;��, �཭�I�P�ĝ�������ԣ���6q�`j$#*I��G��O��T�"�+����ǝ�(5G�.���Ř�������l�S�㫸����}�s�����_}��N�����UV��I;�u�[޳�4�z|e���u�Pπ >�ig���욬���ںo��� ��d���
�x}����S	g��|����l��|J�5��%l=b�ɉ�u^��u���x4l��(g�k�Av�9n����i��z�����Hxm�`�;�����K��ݠ�&㤚{K��Wl��͛YH�5��M3�X���+7����fmL�8�u��K�� 㽹���y�W�d�+��7�?�E�o��Mfez�F��%�Wtnx�7���x��K;�Ƀ�^�l ��=��1{y���5�>�cIr���ɬ_f��qM��lAj��D!�bQ�JT�'��H :3�AŅ���Q��{Q�ӌ*rn�Җ!�]	W�P�^��̢w��pb�X�,UUP_��[d���?�CsH����x�Mb��t;y�텏{�fg`��#��5�������z�����x�V#���{H_/��Yj��r��Uѡ�.<ZI%&�Ӧ�����'N�����m��ɮ�,,�~���%��Ώ�:�C�3O��n=U���O���]`��{��c������H�U��X�I>uoz�g[8ve�&��@�{��ކ� �[�Ύ�����,}���8�Ù��VH����ye ���(�O� ��܈+�A�#s� >�3���3������e�p�K7���q;�������X��Z��t@v��+i�ݕ�}�A����m�H���we�yDg{v=���.��x��"�AA�"�")��gyN�t�F]{��x;�ߏ��έ=�=�V6Ij	d�W�/��cK�w:��5���I��>�ɭ�Hm���7�b����5��v�6*��g��A���u�!6�*�sA��K�4�'_�}��K�����C~>��dQ��y�	��P4v3?y�8^�1��M[�cqp$���&����1�;�q��\l��ۤz�2<�;)�^��&��<c˵ٰ� ��nxݷ��`�.st]�]��,����~}Ǐw��� ����':���&R���K1j�Jj�y�>ϒ�3�L���aA�6� ���n[�ř��8��y�^�&��9�<X��d{o��UX9�f��	P��"�V���-I͝�j���-,��3��JO0��VꩧE.>'�֘q��}٠
���l�=�������_N���Q>�fM�j������Cm�D�XJ�2!�DX
�>��ۏ{�c ��w��ƫy�V���H,���`&f�?|ٔ�7C�d3í[Л�6�����g[>�p���i1#��H䖱�[��\ӚP��d����Q�(/N��Y�? ��fRv�� �6�4����!�p!+���X	��v+%�k_i�<KO?wq���/����gN������ޜR8�[�z�y���}�o���>>��Kg5�{<D0�U������
���]�ƙcY���f�m���G|���jF��WG��������4�2ƒ�1�骝�;���f��@���B^���7z�7�)��9ӝBr��U��x4�
���Oۻ�;�v��W;ǭM����郪[q9�}�$��<��'{����@�ŽQ�� ۣ{�s9��d�U���{����C�"8�w��&��J �������a��o����0�nd��Zd�\��;N�<8�٪f��=�S�F��ש���@��{�UV�g���sR�, I�'¥Ċ	8�b(M���O,2`�yg��y���Rn޶^�r�_E7�xQnKɂ$e�-�~�����B�����o6�v.�Jy�;A�����\��۹21c��RH��c=O�)���9G��`�3}��Bʍ�Fz�1��J��z{2~�б�A	�8�̻���8N�����<{�Ӿ޹"���(,�<���^���G���$,�!�r�W�y�a�~	﯁D� 
vY�l�T>��"�����7˛Ś��XU9��#�=̋0~�N��O-�����f<���<�� #���HUAT7>�j�1tTp�������ûl�6'G��
���8w�N�ɬ�"a�~�fا>���+lUU�"0>�_K���~o8��sK�+�O$��M�7�u��c���v�r���f�tޔ+���菵�d$4�wp}=���TyǮ�& M;�3߳�A@1Mw�΍4߽��Y܃N{M>��3��A {��3� w�<xzɄ\�P� ��/Vb�����oNpkU��β=�%'-w��h��o���z���H��Aj�MR�R��ob��C{b���M.��<������+g�A��D���-�&nvN�WlؗD��k0n]kUˣUGQ�*H�S�9�~�EK�FAv6�t��,Q��-��'�~f/t�,\�\������߃ =Ky�����=�av)ϻ��`���*5\�8M� �&�B���}���t.��[��|"�R�\lv�������g�p����w�\Re@���y3<��n����J��oT͜��bsqRw�"��f��s�+/�W�{�κg4�qЈ�P�	����� �vh[ZRo[>�c�=<ً����1ܫ�|@���c��8�������|���@�ҭ���`�حR�$��8���[���N+��pZٿh����~�]���4Q䟛�~Gk���󩝭7���9C�)T������柹 �0U�)%��{��#98	�|���t��>o������w��l�C�e��rh��P�(l��2
��V���]Z�u���٤�`�9M�j����7ˋ3��&N������[�����_�	�{��Ś�gR������i������rO��2�h�z��9���}��t0YI
�"����{���!�'J'��;����|>�<3%�ш�:��a���1v]�jS���|�#�\|�N���?}�<,��7�� zs�a@F���K>��$���OlM�G�zٴ����}�T3^�o���A���釨#l���s+C{�!�g���dV�_�^�~��ϓ�����*�9$���\9ݻrNٹ�=�uk�sm���bT��Msa��Y�l��j(S��R;lk�c�Q��\xB�zM�6�o%dX�*!8fh�w�эr��5[m�?�Y�Q�I��ܓ��~,k(�s���{�G��bHג?��6�d�}��fqv�j�B�Cߵ�^�~��׆X��Ղ�^Cz���k0�\�I���'�b�D=}#�6��/;�<R؜.�29U�U{��H]!��7�|� �����8�I��{4y�<揜��v�ݭҥQ#/�[���Iÿfg�����@�*1�Ę�oz�ݾA��K��.��� �>�����I|q}c!��|=��u�AP������5q�X��_,�v���ep�\kԵ�T)!����dA�:�7TFg�*������#����0�_* ����m�G��>�;޳��W����M��X����������Zm�;߮��� ��'�u#x��Ó�۟b�6vB��ޫ���$fF�[@��J�IQ����t@�B��{�s�Ͼb���D��=>��s�Q�|w��|��>���"d���w��1j�/��q���?ٰ�[yzWa��E���� Q���0</Zd�7��o�����_/��$E
��7b��]Aim���Ͼ�x��,����̆M����8KM�S}��͞��TB�,+�� ��9���6�k��/���d�"�K�C��3k���,��l3�f���1в�q(��.�ˀ�ރ���^����$���9�q?\s��_g�L�W��a5�Fr"���X3��w�v�?=L��y���K��F��=.�9Q3������:���B�4ZsF+9�W�帓�(����3B�g�~�'��/j������NKޒ[���[��4�矼P�vO?V��o�L�ۥK�8	J?<pa���dw��G:��/��?�)���RQf_ �zt�������ջn���*f(Ǡ��Jz��s����={���P�"�8����ߏÐ����C�"���u��xT��<�e�����kv�ݶa͍�hG]�c9�ccGmt\�|�=:ٶ�
�m�<�r���m.1�S�]����ݻoi�ܭ<���]�60^���pm������îݰt[���n�6�)!���v$v�5\��f<�Eb�v�SnĜ:p*<����d��4s<\tm�v��UŶ8ᘻc���aV�w�v	�۠�s�8i5Ƅ/Wn��L��uN�`^"����oN�� �=�Cq�]��E76\��]��݇U=/`�7���ۑ�{(�9+<=���2�:�V<�`X�k�;���g:㡮���uˮۄۧu�퓉�N��k�]��m������-��.���nK�v��v3��ȮQ9Lsh~���ߨ_?����xy|�]d���`c:r�<|G�����J�hI����G���1W��J|t
�ģm'LN��8����d���1�A��&�wF˓�sq�Q�E���yx}I�2�Ap;�Ư�RC��#�|�J�$�*�0�xf�����KǾ���E�^	ĂN�h��J�!z�~&���?Nx�wʗ�M��u�T�.�6	�e$��I��ԗ>���BJ�{f6@83�� �q䠣�a{�IC`	�6�ї���0sk�j�䱋��(��t񛠑�y^�]���K�V7������a;ű�C��j^5fhN��!E��
�ԩ�����2��Ru�d%M:AA19�A��o����U�)=ϐ���QA@��~�g��K�8���G���}ި;��@�x�3��A����>�_L*����=��Y:�Կ!��T�.׌�qOL`.��أ|��7���flu�E�TM��O���O���x�/�����>���=jS$���jR�`�,ee�T{�ۤ�~����O�zU�;��Q9b����m��_���s܆����4���徜�Kժ��R�1�]�TڈR:K�?�%ܝ��%O~���W�{�>�W�|.~��_+�ˮ�f��Q��9W��zj��:%�u�Vfx�O;�O�w�)��ֈ���[lPI%�Zٌ��� ,3I���7�ςlH��xLG �$k�_y�Ͷ�`�u�U��B�ʤ�|윦;t$�qAP����M��]|.��jJH�l�7�� ��I��W�\�K{����Sf�oY��Dz	���������!�Fڠ����Z����r�39���L3:�Ĩ}��+��H�V[U�X+�R�s�u�V�3��Kdu�N�dI�<��T�Kw���X�|�>�p�Cw���l��Q���눻l�7a**gñ�*��G>n �YȎ;���V`�ɻ��z����K�FR*�<v���	�1)�a��݀�۲��Iݮ�ޯV;{-8�+��j�������X,��vr/�DɗX�u;7NB�a/(�Ds�.�}mIkR�Ŋ��eް�g�<��a���w��
���2VF���m{�a)�U]�|�P�C7��Nr�!�g��A@��G|�3﷢��d���؉�������+�M�6| ��-�6���e�B2V8e��)!Qb���rt^���C��xq=��
�ڧ�K8���SS�y�ے=Q32IH'�EH�͜�dϾN3�guD��Y�Z�{�yHiM�t2h����ag�D�]Tw�߄�#���l�����aa2mh�[U4�2�c�;#���L�x�e�LUv7�*�d�yC�?u�n�s�C��k�c��4%f��z�0dU�9�s����zk��*��Dc+)~�N[;v=���|��ҫ�ឿ%z�S[39�~�SF�8�����h���"hn��)c��:F��ي|���|��ugƨ���P��e�	�gy�K �9��"�zH́�4QiU�Y����{G��ەjA�#�m�1|?~�	z:�v;�*�<3�mol�ɼ��^�;j@A�%n5KA
>!0����i�����΍�-FQ7�'R��K��=��6�{�7c�܅;�39��"eo*�J��$��W�2r�2��l?3 �����6��X����m�*����ޣ�r���=!aKB��v�R UZ�r�&6�PmЖW�v�v�r8^����wj�'`���IBV�6ێ��������DIlL2I-n&�<� �ǃBm6�6�kokv���)Q�@�"�[Aem�ٯ�+�$���N�B��`$d�]|߼�;�G����>�n�g���J��,n���B|{|�]k���/��M'h�u�@���[�)BT�gz���2닧Uj��W���:.0y�wN�(�+��Γ^o�9���g�yDb��KȰG��y�Y��&��j�����&���˻�%���X}�6�>�ظt�l��7j�9M���>���YA� �AؙF�u܃�+_9�|<̛Яt>%�l����y�Jү���t/Q���2�����,Tn���	�D��5~��gf�;|NYl��������z���6��t��L<��>
�8�EfE���K�xk]�O.;��6y8�Qi�ǋ��t\�=jw#@�OmTe'b�}}�?0���3v#������W?X��߻=��p~���~���Ql��r����,K���]]�?�N?����gj2zI�[��?�9��2Q3�VJ6���!�u��hK9��>CˇVÜ��Q���E}�"of����k+G����k����U�0���Yv]M�i7�O1e�h���"=�x K5��ɤBJ���F,�ځ(^�gG�+��<q:r��
�Lf��~~D�RRZ�1�V��s��NԠ�#��f��5�Z�Rt?=�%|dHQ���� 2��;PCe}�%qB���/es�$]�Y�g��4�gAe^�_��=ã��{�ij�i�/�9E	� 3	�z4D�X�=�6��p�g��g�I}�`�5@�͆aYr>�Z�����WA��J��ш\G]�N�\L�+5�>�Y���,��
ъ��
�1�i����H�7͹�$��%����&�֕ū	�(�Q������{#&���dU�k���`��P�IIf���=TyuG{~�|�?H*@Ǹ!�ْ�,�f��x>h�g�sd"����w����F+HS������0������
.\�V����J��-�2��N���=��3�_c��F���π��y ?��b>.qmK��8��_������>F9�y�_�2F��O�7��k����ү���^�&�x��H��@���x��q��[��Gy!٫�~0d��#�	Qiis2U�яF���o�Ň>�{Oh��\�68��,��[�o=VyѶ샛�s�Uv�gk]T���^*v�qqH��丬w��(ꮝ*5�TE��X�m&�֔�5���Zn+ ���Q����r��x�s��Jz�}� 8t�d�r�j��k'�D��&,�5*9W�e1�y,9�Y�ަ4�c��ב9� �*d�UJ�J܂���	�r�C{~��.�>kR4�E^*�N;%�+�|�݈�Q���~�ܯHz�iZ*�+D*�*�� �(�J�c�ig�B�QN��V>��'
6���|�A��Ku�[�����d,9�^��#ͮ/��K)\���V��1��m�Ed�F���͝ߩL��]����j���ܶx���|!u�C�T(��o�ߪ$r�-s�/�
"�p���^���3���1:�ZP�(������6���zt�8�*��}-����C���5$�!�R�7ᵋ���"e����SLV
\0�-�#CyL��{�H�>g�����*(�6o<GVs�J���}k �,��F�3an*��Q�37U��-�[���_��~����I���_�$�h!m�R����QkU*
D�~�CkRV&f���N��Cf�_o��K#���H��G[dn�Wc~���Z>�IE�^-`n��Y�w��r��Oe��=ɘ^���G�'x&ꅏ�t;����-��#�p�f��*,ƶo���G0MvD�_y裏G���W;�_�<���٩�����NW+W��V(�R���Иn����9^�7k��s�\��^�y�sz̐Y�u˙�u�V귍ԧQ���:,�9�Ģ�~��籃v5,��ѕ��R��b�z�?�{�"�؋F�t�ݞ�-�kdզL��8���sv�2k^
�M盠��_��D�O���.,�6z�C�`Û����d�'a**g��AU(�qy����dx$�����zx�.��0v^�t�����>��"�=�n�qU�Jf�WeBY��]��kr�Mk[:Lo�J�$JⅭZ5`�Z�[�**(v���w��x��H߹�J��F�7��ys�J�>��&L�_=�0�T���}�z#���Ͼ���p�M�d���H*��Gy�qz掿S��'�+8�W���2{�d�|�X��'N��C�o'���F1���SqY��b��F>���^��|%�H�F���b*5�Ա*2��k��S:}�l%=���!T�*	���r7���1Ը�p}�~��CJL�E�2!��6䒫^����z��{'g�t�Wcz>Kؙ4SS�uй?6̞�ϩ��:��3�=�*Z� %�BG������g{�Y�+U��v�>� ���ص��UKcDjV��Q"J��|��Q�i#�S�w�'L�%�}�My�8�m�1�Q�n�UNq��\��߳-�sK��Y!�wV !*>*@]�G���Q�n��TA9��#�z$f��fJ;���^C�{:��4�����o�$�ˆ�)�?��v��u�l�Zuң�����N�h��G�F���yn>�����/��9��H�䯟n}�f8d�x�N��d���Yځ���y�Іc�ȷr�=���A����s}��x���k~���=v/<�r��߹H����q6?�'�T
�/�GW���kg�}W3T�,;'��-���`�~���Y��ul����YA=�9uJ�Tce�g�>�����ۜ�"��z�}�_�Mc����oe�?k�d��{���g��w�zi�^5�8F!������|�������pn5m���lk�$m��⨨��Ӡu�o��:�6�QkѮS�s��5u�u��M����Xr�Z�ɪ;�9-̭u�S�l��{3�J籇����׶��h]V�v�5,�>���ngl����S���q�z��^���^+��[�s&�6�ۮ�sꭃc���ڂ�
0v��d���J������أq���y۳�g�]Y����㫴�le9y����F�봝d�v'�u�\Ob2�ryh�{9����]8�8���h=�G;n:�:�A����',W�@)�Mݮ(� �Eq�
��%�M@�jӷj�@=f=q���J8�k
�5�ܼ��e�Wr:�"[1ݩOJ��oO�砅�}��2�)ŏ"q��dC*�h^���#��p�5I/�í���7]�x��{=8��yZ�I��Z�g{l�#�Bさ�'Wr�צ'�!(8Cdϯ�{7�ӣ�� ������dA�~L���NdA�t��a|�,��2t����!�m�8k	��[F��ȁ���4�8�bzl���xV
���SA�b; ����R��	���n'=�TJ>8Y�1�42���5�<��׆1ˋ�7��2�$�Fv�9��t��;r�=WO'<�eD�ss�@��]�e�k�zbv���i�z������v��5n0��yƴ�b�m���Ŵ�D�)K ���8k���}�Z�
�l�uJ�U2Ek�5�ˢu#�CD�]1B�����H�>'�+8��/��L�+��4�7Uc�Ř���g��>�>2!)'u3�Eƶp�_}�vYA���}rq��;y��;vn�>��n]/@��f���k]z��K�^�Ud[>��r�Y�L;��Q�'��NمF�6������mZ�j�ڵ����~��{����ͯ���k����F��l��K��lɿ���7	P�� �`�R�e`��}c����6�γ���bc��FU	(�|�F���(��k��U
��`
.�n|�t�m�'u3+ʁy�Ǻ��<�9���ċِ�}�g}�6�TFKB�Z��-��ʕ�Z[alD�TR���x�׾�}�ۂ�+~�C�7�߀	^�H��pa#5�>�ѓl���8��P�P�rG��qK-�\�~��xF���8��bi#&���y�K%��p����
�7`.,�6y��6�M���Sd�'y6w�N��銩��y_S\�L��{�n��4���R�F�)b�EZѶ��ҵZ�E�J�c�@�����r97���]���3{��F����(ʜ	S&!`BTOrd�N�l�D�\+�&������7U|�վ��|\/ ;��]�H�S}��Z*����7朮��}�� �Y-�dϴ��Y��y��'�Qf�a�'bws^҂��@��e�`?Q=���su<�݋��e9�@:��/+v�x�ɇ�S�p�G-F��WO��u��p�"��8%;vdNզ�;b���jTID�cc��kj��T��T[e����^��m["x4���R�6�^�o���Y}��}����?R�Ord�����Z���w�-��+�0�i�>%ܙ4SJ@�����Q�o~�y����L�}�VKN�e@����I���ؽn�ݏ�鴂=�>�x�{غ �v7^�y牒Us�ܟ�݌��K8�m8�zSD���4)y�y�=߉�/b 0��Lx4��UH�Z��6TX%/��M���|��y4P�7[3N���e6x_xꩅ^�YC�4���F���B]t=\ݭ��oL��޿c��l��.Z�i8��2ǽ�#R�;�>�3��_2!)&�|2T$|T���wߨ�7�A�ӳ�8�Ƅ�O�Q�~�g�{�O��u��͏g	ЇM��il*���XR�X5�Zت���&�9�3`6d�����=�qj�|���s�ol�ɼ���>�Y(�����lU���#�;#���yM��pgS0��m��8$�G-��]�!y*���˟M���બ ��+͝����͢:*����f��z	eH*(���V�zv7͍7쨏��@$��%��J[X��Q�Y[j�j���ѥ-��|�vL+�Rmag�Qp��FG���K��`5j�	�� R�J�B)n!{�y�K��Bť�:��BD�sτ*(�6o=�����U�٥���Q��>��Fl|���y�K�쨃��Ψ�4M���A��͹��4��^��i������䋋�{��ў�$�d��bT����JNi��Ol�%��0��[�s�lV�����Z�]rgg�Y���4�S��b×��#�V�f��J�F�41����i��0�����ՠ�[m�*�Db�ť�Qe���f������BU	+��+SL�T%I���!+�Gy.e�p \�冀�FD$7��7�Ϙ�1�����k���zk�A�]�-jw�w�w���YVG"�� ��&�㽢p}1����iOKظ�_G�p!wp�GÇOo�75�g��[˜:���jU�2��Q�2%eih����Vڪ�""�Pig��;����Ǟ�u���c�_<U�|!��ʥ��|s�7��k�<Ħ�zz�����ʠ�ct$���0R�sI,v�/�g�bS�6ϼ[�]ݡ�.��k�Xn!"������+����c�2��߄�6�)z��c�BȄ��t%�Fq��{�o�8�w�:�*�{���y�t��O'⻻�<7o��O�>��z�&ћ�6����b��	��Ε�KH�}}�t��H�7p�ݾ��4gu��z������~��N��=��t�����7)�k���'O{�`/=�&'��9��-,G$o�v�rއ��ޓ}��n����:����]��~�x����X{�v#�sg���/RjC�s����7J��㏿;_��s?}�3�&�h��oY�d��(���<on]��$�?M��7�����1��4J��C@T=�_�xG�m���Ӏ�Fё�^\��>��\:1���y�?iu�ڇB��Gr��#m{�=�C]��CV��z*j����Q�w޹^3����Y�9��i��V��RI� #�i�kΝ\�>7T�]�WMŹ�t�7Z�YD��
@Ņ�4��{���]�>ܸhk<���^W#B���u����Ϯ����V=MR�X@�Q3#�0��B@��)�>G|'�l:��>\�#��ڙ�f#V�k��n�@�Ow��ݶ�m�%�X�[mJ�J����m+-�}��34V�jq���nDcd�T#"��M$t�����A�g|�ؾ�+D�9*vEX�V��"�Z�q�7#�^�cg��%���y`��a��ɚ�'�#��2�Q⋗bsz�F&D}�=�A\���f�=�{Ҽlk��<�.����N��<�{���(��UA+Q+Kh¶ V��֪��$���`��{�ﾶ�#�ٯ�����H��
8���%�8j[�+��$_<��Y��z��j����/d2E���w���lϝ�#��l�`�& ���	�I��"�c�}���k��\կ��#�Pv4G\����W�u>�f���������I��H� ��▕���&��g�ɸ�zz��9�,�ݵ���]>kv���`�v�%��6��Ѯ�$�ڭwa�$�m�<�X�%PQAyj�eB��UV
V�Ъ
�[R�[R���	��Q͎T;m��3Д�
V�����阆���>O���|��ݖ����I`t���8}����h����fC����f���t}�%3�4�W�'�su  8J�u����pɃG�٪o� �Kg���Pꉦ1�l,!�Vܲ�\��nL�D@�f���ut��o�y�z�:EU(�h�PAPX��h�%cj � �u��/�}
��5���T7��H>gWRM����Sg��}���&�r��y�2 ����\4[l���($\@b�Jq ��:���־�|��w�}�}�)�S�\�l�_�}�!��b�=�6��w"�/~��a�}�{v<����s2�(�X�,b*+-�EjX��~�����?v����*� d8���K#� �㓴(��\d�R����Un83�9c1���ǎ p��/�%5���1ܶ��G�=D'<x���O�Z޳^%��6 =�Q\�MߗtD���Wk+���#ƫ�t���ͺ�]��,ET*UUUX�TF(��"&��go^��)�Z>�q�f/���l���R	�-l*x��w �,��:i����}W�9�X���~�������*W�9š�z��ӛrt��÷$���ۚ�c���J������5ڞ����cǽ�~��_	����߈ی�|����nb:
��ֵ۞Lڑ6<������j�p�cٻC�ō혮^�����i��e&vj��:�����f�V�x/��FҢ�ڪ�1F0�E���-J�"�k�幻����vl�(:8����������U#}������?{��DO�9W��.�d��
����k�>���u�s5����1{�w�'�`�e.IkF Ը�jj����k��;��_�{��B�4@��_	κ�iL�c)ŗJ����d��H�c,�QBL��$�	 1�1�(���(��{��H�c��ּ��s���}�x�妟]'���܄�|�}>z;�����Z%q�$xm�͖��a3(&	�Ӄ�K����|�tu��$z�W���S����!��[�9�&Rð���(駴����fgY��йy0c} �7���DDE�ATH��E	 �y�:#�ꙅ�x��5P�I�+Nx��4;��U��5}�� �	[����*�(U$ߝ6�{�J|{�M��$w, ϣ���u�U�� |>��FB���ա�� {��q���N=�j�g���71�|�U�����v&h����PUH�X�+	�I �r���aB���Z�y<Q@ux��Ԫˈah
U4:�m�J!W4��n��;E�2���Z�Xh|}=]	A�=i���3S��|!)�;��U����N!H�C>W�1X�(�O�=U_-�n���%�	�>�鸥w�V{VpWm����m:x_=�j�T�-�8u�#{��^���ߊ�N���;.�P��/���or�5��v�\� K���V��#�_��?3۳�EdR�f}o��b"/�Ő���xw;�|�-I��w�l 4��fk�܆G����nDƴ�1{�=�+)�C^�Z*��ܾ����p]o�?M�O%���ǚN�S$~G����%٣��'o���S����s�M�����_^-�	x��zf��<������wi��w��	�g֯S֙Z"�l	c`�kԝ��w8	�{�۬p�gpn���Xs<v�x�𮗨�D���/��Xi�9zuƮ���n�zSm���x�GZ��q�Z�;y���A�6�]Υ�ƴ[m��N��k��nNJl.�w�i�컄���=<��ٹ5��qd�zk�S�{]|83�Pc4�q��ݤK��Ӟ͞�v��Y<ۓ�\�5[cĖ��^N�!�9����h�Wq���ɷg�cB]�픞ϓ���۞�6KoQF��=b�,�r�<
`j��۟��������̃uE�<Qv�֦]�e�.��$�۔���CH푎S�M����۝�b�t�<�Z�a��Q����&�t�ԋR��]�e�	�cd��evc?Q��y;��W���@}$���aS��cfam�&R!�}��~>x2�ĕ�%���)�W��u��0������P�y�ؖz]��^�g;=�c��5�.�sc�O���p��Qh�e%��ɣ�&� �<�� �`��c.PAcy2�gm��J����G���n�uz����;���:�Sܳ���)n�q�f�@~Q�MW�3��7]�kʱj(�Ś^]K+܈L���pc&���, 2���R�G���Ws��5�Q܃�j�:����WR9:��On�$v�n�m����0mS�݊�{qx�zP�\b�U(��a{k�d8U��F�È�V���c��KkZC�*�e	Rj���5*n��nJ���ƾ����ǿe�����2~�p��Fx����O��'6 �(����uQ0F�τy�,"��w��� 8���,NBG,���FR�5\d��U����ӟr����x�F ��r!�7ᱦ�O�j�ތ�je{Ȩ�*����͗�<��ofo���X�Nu�S��X.W��^#�KB}�����'Z��>�/;9eq�$L��(��V�q�J��׶��'��m�u;�6>4_+3�}���do/�
�4���g �Wn�E�n6M�^��i"���mM��&O�	�I$5,�D:���&������_|sT]Z| Ϲ`�e��|k5�|�`�¶� WF���q�) ���D��G�g�-oa���'�t�p��.�!g�������M��{ύ��]^%��:zz����6��oF���V�7���D�I �~6�&�&�՛���u}N�I-���,p�adL�JR�Z���v{��ֻ��3�w�|�p�� w'�����)7�ǹl��J�V��ڸ����r�+�[f���V�}��i����-�{�r����i����;���暌��I�0J17���㝎:�vy�e:�v��8�ͳ�#B[>��B���%�Ԗ�W�Ԩn0��ls��\��.٩c[��w}����~��3����׃	0�v�+�_���G�#5� �dt���u����^��Ҡ��$p����Vs��Tu��S�V-?^)��4tN��f4�F��*�|g�>�#g���Dħ.�V�����b򕍝�����d��>���)?��t ʳ8Kps[�sôŞp����v�xw�$f��%}ܰ��h�>	�J*�
1��ʭU24�PM���ؿ����(�����GǤ�a�;i�^�o0��*LS4;}X�ʕ�U$��P}fǱX��DH&;�
�N�^��/ܫ�I�䕩�����j~ϻ�S�
aN"n�
7��ㄩ�_;	Ňuw�����.﩮]f)�G�(fl��ޫ;��R��\;
���21 O�|-�=��ѷ�^h[��[w{_^���>#ݕ�xp���������Z]�6�N��&�TU2�5Tp��Jm�t��Z��o���� |>�-��5]f" Ο�{���ݳ\Kpf� �)���/�l��$�����.�W���=��
*�OS��X�#�vԭ���A���^̟��V7�<X���	�lޖ�]�J�{-:I�O�짳�7���Jd˞c���ݳs��X�9���fn\�k��{�=�t[�:p�����m����JG�`�������W$��R�L�zir?Ew���t������H���]g�V�ܳ�C�l,���@�� �E(ʜ	SM�� �s:�;��ܥ�J��wt�;��*ǎ���!�[#J���|�J�q��¢�C�A=mE�<I��Tr���{zO:Pπ�OtM��]��{�,�>דX����dM�Ȃ�"G���=�]������z�ލ܉���V�A�ST/�K!�WH�ߢ����3��=�NBC���MRD^�|��~�wp7'hx9o{���������8���8}��R����r����H�ݗ�����I���-w��ct:"઻�;�9QDZיX�r&ys�i��콏_g��{`�H�-��Co]j����>�O���F����3�{�}<�[���o&Y��lʁ�vK>Ǹ�T����@�����v�� W��H�HCW2f�7;Kg%r�_C{�S������d��_����9j]\��y���{�嚰�����k�KcV�d�KQ a�)�����9�z�&b����ؼ�d�:�C���U��6�v� �r��:|�\�ǫ���gWk�2�՛�O�{teh��w
\���;�_�^�FE)ْ���鲣�ʄs<H�DaY�!�7;fy���U䘙Fm�E4�<�bើY��3��N�E�ӣ���]�mͥf�Ք��X9�3�0^߃Av�m�л�`�Su�#�}���*�y�|�m<�]����|g�W&�����ЕT Av�ǪD48���;��VKpc� ���g���V�݆\e��6(�j���m��Ӌ9Έ���ڰ'�z�P>&x.vЪ�R�\:ib�o�z���(�Q}3�����z�h]�G��aF���	 �B��=e[Nvց�cH�S�����@��˖�F�����Dߝ5N��=��<����q�5j~�:��I��U*��,Y�����j�Y
~�ݭ�v���,�b�$��cGB���ޤcL���8�H��WX��h�i�喐�+]u���ۙ�\�p�en:�N�T�]M[�����gI� ��퀹��&+8�������1q��v�r�\=����?\�=/[�N�H
[,�;t��)��[��<�'�y�$�������P����
�jw�X��*���"lz�P�^iϫ�D5#�π�z_���uZ脂1�H�,ce,��0@�nJ��zkGF0�9�`���\���8b�DǦ�G���L뭣�S~�qy{�	 �s�'���x��$du�F��a\Lp���e��-�@d�^X����J9]�uw����
�6�PYZ��Z�l�i��CN|�Q㼆"�ܳ�;�� �'��X܎"!��v����5S��	�5
pI��t(�����d̟� ��AZ�f�"S���]
�6G�P�M|��Ws��f_��<Bv�VHD��7�:9\�}�\k�ܞ��{�I�'<�|}kid*�zǑ�4H�^6:]�=]D9���COH����^���й��y^�N�n�b%{��`xH �X�jރz�����ePw���m��w2r�䶳�J��7C��[c�3+w��r;� �fG�͓�I�5��=kDq�D$f��Fr�(�(.��<���id/}��c^?.���켻�Oզ�L͘ܓy�;�9:�h�5۠�ۧ�v�u�r��eפ��o:Űn��J,�ۜ�透;�l/;�w[:	8��n�c����^]�q@�::�������q����UqG��Y��SLRB��o�O��r����ӝ���P�2'����sآ�r�W�$���><D��?r���w- ��RG��o�!��f!EkLNR�m0������T����!����3�I�1�Q�)�)�-\,��V�rz��V*��;C�'�Gä�
�,ڧ�6g�#�P]E��Ф}�T�t�|��� e�S�bt��E$��A��Fc�����NB����)������W�W���,'
Gr�F(h�[ׯ�Qf]:���e�Ӿ57���$Ēf8%��$Ͼ�5�,����<v�3�Y������gz��p'� P*�	F���F�Ъ[9�y+�W�)dm�qJy\*��è�-8�T}��H�N������|�Hw)���z���#�����6�0m�̭���eK��~ �-u��`5E��`�\4�,&K�4aj]M��l�k�z;��"mq^������ϖJ�9�Iu��'����Qk���L9��[���}�GX��	$}��ɿ5�̧�G�����?����UVHA� "�P|��"���4�P��k������O�ܭv`��Z E	 D#	@Y0�P�X�Y�B@j �EA� �V@Y	�T�@�@����� �L$Ad H+ @@l�T�X`RR� u���Ao RDPAD$A@T��E$DE�K�ʨ�x�Ij#�Q�Q�A��r�2 �h�����$a@h��
!h ��^(��@"��@R�@
�H2�($��Jyጠ�`n�X��M��G�PVAq�F�O�����m2��g�w����o���|q�}����C����a��ӣ��{u{�pf9����{>.�U�99��z~N�^�z��0�F9�9? |?�O}{��D@E5���=����:�=��v!@{_��x�yą�u��S�T�'�u�����=����j`�C�d>�L(��g��	T��e�2�#�w��)G(��u�b��� ����$��$ ��D ��H�E")����@�D�A"��0X(F"�R� �
�`) ) 	"�H# ) 	 
AB(�����Pb� AR ��0�H �I"�A�"�F���	` �!I@d�D�2F � �" �"��
 �!@`��@� � �`"��!
��0 �	�A `� �H�P��H�P!HD�`DB �A����� A�@�0"�+ ��`D�� � �*��,b�"0" @�H� �0A`�0A"�DaH�"	"�$	��`DR$ `D@� H ��HA� � a" � � �$�!`1�A� 2 �1�A�1PdAb`��H� � �H �DA ���F
����(�d���H� � �(
 H�F�� D Όx-����cu�`g3��1��?��z���� F_!���/�j�����N�3�j=�C̝)������жռ��* �X�!d����G�A�.�$�{�	g~FB���8y���,�GwRk��|�/hj�"�r�#x�􁸞��x��5��x� KΧ�PS���F/���h�V��p�����p��7C�J��ء�`_kPE5������=A��g:٦R���� �xL�C��
5�8T��l��ǿ��;:y� �v����t!�z�R�^���?_���͂�#q|ު�{��|���y����yߝ�4���G�0�w���� E9 G���t�jm��'��u�#A�����%�cGY��r#�w��n�N����7�-f��T��7���QTs�o`����l�p46���dP<	��7oV7��#x1DS���GB�w8t;�]� @E9�[� ��ǵ���þ9��s��\A�v��_,	����nA?����O����rE8P���%�