BZh91AY&SYQ;��<�߀py����������`�_��            �| J(PJ
 �` (( �à}          	�  ����v{�{y-4�Ow��s:�ۗ`�)p�i�oq�;� �C#&������v�
�G�� w(<��dŖ�w*��Ϋ֪��V�e׻�"$��ִxn�15����4h�&Z<�  ������&ڍ�8nr���\�hxwr����Nܙ��srY4j�և�u�\M4fjx
o  �{�dœF6��I�L�5�ìSNG�T���;���=y�ƞc6�ì�΍h��9D��@=�wx��k�s�-4֞�㷏^t�^I ;�6��r�Ow8���^��U
|�          O J�4�CCL�i�Mhщ�i�)�`����Lh     L  ��RQ�` L� ���"{J�J��z�    4   �IJ	����0h`0F�
J��0 F��)�z������S��y�wׇ������˯��?���H�����$��/�X��������/�u?�����G]&����wN8�'�̐��j�X��N$D��aُ���i����D�ܩ���������_��	��g������ż������@�˴����8����DRu���5�^���vq��d	;4d�hw�`tPx�@u��XY�}v�$\�K*0vƗgjǽ�^�[����ƾ��8d&�����V��e6
V����&�á�r�+^�d���w�W.o{R�/(Wc�H:5������	�5�:W^�NS��dΜ���}��w8G��Z��]3j�;�Y��yw�{u��ni��u��f��ӱ3B�C~�Y��f�qD��h�.�����vǫ�,L���0]ǁ6�)��:�a�΁[���F�V��O��'���y>}#�����Z�	m2�=+�nh�!!�OSBO&u;������� m�Ю��ƇɜL#Ŝ���8vi��U듄Z��goQ�s6j�z3�g3��0��R.��թ���v`�&s=;��b\��u��������z��;(��#�zb��Z&왧Tcr��E�%
8�u�;P��9`V�[ ��u�d6[���9�����tWH`aظ#���)ooN9�p;��Ĳ��ݠ.iv廷��X��1�(ҙ����6�q^�BZEb|��v2��G��?�#���o��W�8�@�(7�,�u�\�|��P�Ɉ0h�d���1�s���:W�����&vt:����łf�nn����UDT��Y�B�����qgE�sx����B�1XVv� ��wCKg��I�kf,F�p%c�*�t�&��=[�vs��vs���M�U�gB��\]�k��K{��P��I�`֯2�zÃN3)��[�Ʊd!pقjV�}3gCb���0�����\1sN��J&��h�^$�:gv�}�;9�� �)�_EfWr�ke\����3���s;C�9��jeAM$vv��{q��^qzsn�=����J)�۰��F��u����+N�:ghƟʨ��d�PGaӚ��h�O�����bk�|�_,=�݃Tz��6���G6���ɰt-�[�7��)�ם�4 d�&G}�/p�����!��m7�r�TE�vm�˨>��|bA�I�r��,�J�N��U��;���0s��ë1��ܺ�����61^Țnwo���øΏ~�7�/��3��Ƣ���9Zoa��<�x�5��u�P���̴�{)�<Y�%�.p�:I�#{�K����u�L.^�����4UA���I���ܿN������G��Qr�6��4J�l͛��DC��
%<����g�η���C��N��xi����@�'9�\`�Z�qJz���8�q�Cw��s۪�n�<�Ѱ�n3����uSN�A�����dŶ.�1�Գ���6���'����n�]/v΁MbvE���X�+�L�ٝR;�������.		ݢ�|C;�ɞT��o=�w��&% ;z���k�F� ��"s!a�����l��5iʙG�Y_ ؊\�n�\�u��7'˙FЮ�O�j��mL�VT��Ul����kK$�Τ�(�CY�!N�4}N٣��.9C1�o.Ǆ����*�'���4��l�inj\���6d�;�@w
�1�%����e�a{4��m��7q�����u��ˆ�q��۴Ǯ��s&�<7��R<�x�<N[�.��:�فb�N��4P���8��ݠ����m�Y7eSg�����c�t6�*��C�.]}��[�v��P���q}��t���� � ufJG\���z��E3����v�Ӓ����v�E��>|k,����W$�QK�%�4�9"�o$MN�����v�+5v(V��,��LHiGT����kvP�on�n��ܝa>�"�)��~Vq�f[�C���\�>`;OF����w����M$�:w 90����:l����V�Fqqp���uK�B�qm��Í�ld�ӫ�g�j��g@���f��#X��͒���3�: ��"w ���NL�S�$< e�Fn��r���i\0b�"�Z�F��V�Ȍu�9Q�9��Z_i�;`#WJ�K��o�h�Y�A��ph&v�û �ˢG*1eg��+e�u�5&���ɡ�ع�+�{O$��A��%k�]skvJ�R��]�c�:�\������0��\��2�r<aH�)m�Ŕ �`O��;��d؝�]O7W�i��*�E�ب�$�9'ݸ�Ⱥr�1&�<��{WZ��U�^/I���@8�BZN�g;�4�T�'�{�C�\�4C�	q�7�;{+��  �6?��8��L�دX1�u��J�X����A	�A�un�s�ӭ$��t��_=e���Ċp�4�>�S�N{�v���=��ȕ��k[�W�'�;5e;��,##0���w�������_����n7���5�k�ǰrv;����W��{ǳ՜k����Y_��!}��Y���v�V5F�%kb��R����"��;LpE�s�Tэ�b�'<wvݲ�8��zͷ=�l;�x�:o20���Sz[���S��q,�p���l\X1V�ʶ,�h8)U-���nq]��ݳiQv0�8��{n��I�2�ծ�C��D�H�h6���q�]�۵l��� t��}�y�x��A��n��nۮ�q�qw(t�ѓq�x�ܜ���n��O���~_�������v�z�9jޮ��sqʝ��ۃ�p���Y��b�Gn,ohڵ㮗�;<���蝯�{��݋�3�`�Xқc3�(L�Q[	�:%�$k��97�sk;a�u]�k�ט/�Q��j�C��=�'���"���|�1n��涗k��mɃ�g��{_}����':�un��ub����kkq*P�F[榲����Uq7S`�-sI�E/�d�>�ؗ��n�m��=ex�r�%�<���J�G\`�QF�V�bΤO1i�y����e�66�b!ݕ1Ńn�������x�Vy��qq�y�Im��ۏV�q�۪��L��SS5�=2�feN�U���i�t�o��;���7B$;k+q�o�}h� �V�6���^m?��}��69�l�j���K�֍�\f��U�?|]jM&Q�2�
�[U�������9�]��Qہ8��g�Ӂ�3H
��d^q�>N`n�ց��~3mg�� �d�nzxˮ��?�G�O�v�m��ct;�C�YG�vO����\��vg���lZ7a���u�b�����k���.��Y@.�v��;4��p��7�;wZ�?lnw�!*��reJ��%\q��	l��w/�=v�#h@ !4!F��0�&�":Uw ���=q85��ro1��;�9��>�=�ԇ �`W�49s����xyaU�$����ʝ^�[�WX������.����'h��������o:q�Fcq�V���v�N�B&��V�����:X�-H��N�X��������slR�8^���x�-�72v�]f���fy������.l�����]\m�]�L^{s=yy��\n�6O�\\P�qƣf���fcr�:ۻ.�7�mpxJ�g;�Vt��][����ͳ�0A=�ܵ��Z۶��\��ۘ�������T����;��pI�\ޝl����uLi�j�宑2�,v
1�K~�s�zNh��r���/a-�nw���Y�x�m86Nm�9M�.λ,ue���Ǌ.^�������������P�@�.��ҫ�ɱlSa㷨��'Nq���s���n��q��z�t������܍�v��X����<�97�wQ��V��a.���j�n/:}Ur��+�����8�p;����/��N$��ݲ�c���Q�:�o/k��E�p�sӸ��� �K/V".8M�v��(gm�Fß])����nJ�|i�:�U*��fUY Pቌ��E)+��O��!��幎�;;�.s��ʼ�޸m��׏c6z�)nyez���G��-�8xv���ڃ����MOv��t�z�Z'S�"�RXV��y�v<���9z��:����0��Z��ܗO]�ź���'��f�Ol��[�o;q�!��\n���b|���p�S�Ӎױ�!�7Gm��qu�O�������ܙgg����*~v�
�m��[�����x�w�t�����5�y���`鸲�n�t�۝�#-�֮�n	� �ex뮲���z����;��^���>|��8�{l}�Ng�N\�Q&����gJ'��t��q�?����������㟧�.���<�~��L���G�^�_ Ǘk���{,|63������o2��oP�x��������)i�]v!P���E�������x���E���Y��uoyR+�m�������]�G��gv����9��<�u�E�׫��o�^�
4��n��,fx������a�no��[=�=���g�� xc�NU"^���~q�������ROi�5�����M��T:n==���{�5�#�y�<�ý��'�9�ӜѴ)JP��[ϐ�p���n.e��ν�u�u����c�G-�_�x=�=k��P��"}��Ys�m+vb��!�Q���{|=�7���M>��>գۯW4�u�&ｏ/����� ��xKKާ���~�yP�,�f�p4������뻞��N�A9v����{\��;x\�sO-���x���\}�wZ�Oz��8�k�U��{�&��-�{�����A8�'��mZ�Z���^]}��i𻥞ݡkN����;\�`߽�L(j=�/����s�G��w����b�d�^;���/�^����y��=��NV��h����ܷsr��x;�ߪ��.����#���	�{}��r��.�[����͒��C��`������NH}�o���jg�$�_wS�V������1�ڣ�:_s#�_p�I�b�H�&Ż�I~��A��[x�>����0�q�Iws���eiѹ�r@�'��!]v�����w�������I��\1p�b�׹���/�����=��=#Q�N�Ђ��f�yۿr�8��������K��2�}��tx"{��9���1(�z{5���u�����:��n��<$t�P�7��f�<���|t�|=S�C���k4i�E��n�������(��o����������oC��v�%t	�FS%0RX I�ˠ�ʄ��'�m�0-�=�>xO��o���%��4��|��ɉ.:]���v�Y݁�ddc���$��:\���{y?���7���Ȳ�f�w
9�-�����<u��G�޳��{D���7`�b�g׼��9=J��wJ�[,�K�Ow�|ħ�|<��y��|Wv1����Ӻ��A5ﯻ�u������[��4F9{�vo�z(�,W˃�>�W���y�U�Tz��Q-(��8D���&�FG��}0{+���/nw�fƢ�wo������;��KC|=���_1��=�Y��$+�^	^w�*qw0_�oi��*|�̎��r�⎬���pZ�ৗ������d!���]����M;�v+7�b�}����4m����O�^� �R?g���|ƃ2��{�g�&~7�ym�٪�R�w凳s����f�3���o����Yڟ!��v�U��w���8e�h{����C�Oq��Y��t��[��oz}�Y'{4~�p�/;�һ�wwsgp�,9m{��J�g�p[�	ٸ��/w{�jc&-�����hZ��Ta)��W���Ɯ>/��*�Hn��	�ك7��\�p�i���d��n���o5�E;E��<��f�Y���n����S3ޓ'�+���h>g��mǺ7]��z�ۓ�����K���=�� f����0)ئ�j9�����u�K�V�
�}��\MGY^�/!=��j��qqb��|@��+*�ϲ��x{��[}z���M��s�*������Խ�wH>��,O�4���������d��ўgΓ�W�Ӆᾘz�rۗ ,���o�U���Ro���oQW�v���7qMy79�{��{�7�>O�[�P�<W���}[C>�ȱ��g�}2!Oc�)���p%��F�R=`z`�	�5L�!�1���A��!{9�񛸽��'��']X)�$"��yݠy�w��{�:ǅ��S�=G��+34R<�Ѭ�<������{�m�x��,�����^��z��3��{y��qvz��N�o�_w �;�/d[VC�<�> >Uˠ�ٻ�=�ν�J&x���swoP�h�mζ��v�{��x1��~���B{�Ồpk��c��W�YH��s���t�3f�뛶C4L``�<���ѝ��B�w�='/5)�gA����3w�q.u������ܞ1w�!p<z�e�ϻQ��%�E��0{��Ԏ�L���L�tD�������<1Ѽ�9�n��!1���ω�ns��[��\�/�Yݾ����^�<=���r�&�N�V���|�Puz���͞_�����fe�����Ч�����7��{�X-���zŌ���y8����=�*p��dJy0%*s�*�1�;C�!efe)�V��
��C���*P9��g�� >�� ��ߗ����s��:�����c�ϣo���}���/��>���la��Ks{r��"H�j��S�d4��M<P��j�
�K�6$���^͜��㱒�luu�78��u�bq�_v�&�.qڎ�Yы�]V�sɼ�c��b�&۱�%�mcl�mnz[VW�;:y��s�n��8 ��ە�x���Fٳa���ӊ8CFxG[��8�%vҘ����Z�M��}�tY.�s�cڞ��(`̻�^� ��g˷��OH���tl�wWn���^�7l�t���Uc�u����ƹ7c3�ک�.�깗cȻ��ש��A��]�qZY���X��s�b�T2�P5���ݶ��3\�.���Q����R@��}�����{���N9W�1�f��X1��\{��Mc"�x�K��Wܧ����V�x?]U�{Y�������C%��MH�a{��.Z�q�W.��ݟ���ڡ��X={}/1�[�=y�����h�x�� �,x�*�v*5�� 9��Y��tĉ/q,^�ta��k�Fn�̌�k|<���.:Ş]��7T]S����M곗b*���{�y�F+X�6E=kl���:����C���x���#C|��=�_e����ƌ��d�﷟��2���*Ft=�s�1+��/h�Ah�3���G&�m�svϚ7O�բA6_ �����Dv���m��TFZTA6C{�̘fa��csZԵگ��[3��$|�y�tz�R���W�?u��z7��s�ۻI����� ���fL�o�.[� '�q�&�m��T�l�`Ѐ��k�P}�a�e�V�HD��.�3Nn�m�.�]���K�V�ֺX�a�J'ȢX��R���/Aߞ�/Z�;��wL�u�x�
B)an�F�����h��9;���(�r1�im�(��<Rs�=q�ev=q}�r�	�["so�s~5�:��^j�iӴ��}}t�OFx���'i���c*(t��k|��Sl�1��y��{Hc�'��l<<A��(�T-�{��Ůa,�@�h>� R��V�-�Ǧ���N�}HȊ����2QR!��˶R��1�Y\����Ɩs%	.ݲ�Jvj�ˬ�ۄi]I�h�6m��t�3;�9����m�wlDc"��U��o�f��{y�6�G�ЮJ�au���No����~}�^�����/a� -�R8�Ex0s�6��@XC��d��I�d��C���K��ѳE�O�`ӟ��gs~�m}1��C��r����)ݳ�N��Aڶ8��q��od�<nu�s�UVw&V�O�hoS>���<.R���w0R(� �)����B�0�2� �-��.��ww���0��.p�O�g`b�55�V|�Mh�1;��5K`�]��a"c�L�\Gw;H�qUD䴄�Z:F�o�kr�����w�U���Kh��gUp����Z�<��y��e�\�p�ohybA���k/̬�G����P(�*����g.(�xCuP��Z��цǪ2�#��:P.ƋAPp�)�R+]��]�U���nO�#U�gx�Q	�
����tu�6�S鋲� ��z�4�ۭ6���f��b���UF+\�{=�����M��A�x[�m����W�a5!�����6z��i4��
/S��E�a<%\����m,xa��@�aQ�x��z�e���u�>��N���_������xaw����;�ۇcࢠ��m+V�S|7���1m浬s�[
��%�K  pDtel;���[�F�~l3��-o�[G��`1�]��#Y�6#\����s� �Ǎg;5�3��A�7��rĻ6^�����;��ur���3<�2�'ٸ�)p25V���4a�!�z�(ܼ)�s��y�nI�Bڎ�a��c�8����㯷S7�t��ZKSU�DTb"���6�[o6#y�[�Z�Y��)HEAZ:[[������y�ݽ�HE��b���{zI�]岆z�m.��S�:�h�1/�轂��"1�Ü˝�۵c�V�2ւ�Z�S;�.�#U�^��JBw��A�93e�C�_���9�Q���	�q�� ���tQ�Z��]o�ۭ���u���uu
(K��(�"���;Pٷ��Vy��_n->�w��@�W-h�� �TB���żcq�}���`���O;�%\��d��K��</�����������ƽ����MR���4X�f�%�r�����Z��[vx`�~	m^1�V]W/����Dt~�G-~6~�5�5� �v�.C{O=��1�}���[���Ȧ�T��1�"�	�pѦ�m7���#�7�e�M�۝�y�]�&9��"{��wޞ��܄�%Q�-��׼������@Ms.���t��b�_���{�����aհ�Εf��i{om���/��>ҳ^��7Ձޤv�G�g��0�ysѠ��}(w��N�����D>�1Pʺr	�w�pVv�סe��Lā�'B�v^��N=t��/@{���ٕ{e㜩~�m� ��v�Y�_*�Z}�����ϖ�o�t�9,��.���-���l���s�ѓ޽�Wx�Y�_q�w��n��o4�^h���܄�#��a؈,�m�,2ҁ��yL&V����a�A g��''uX��Y��@Յ3���)��|�Q}��q�+�.��b�DPc%��0�)��,X`<e��,�f+��}��h�Uc+Kh5�V%OeӍ��dPO#���[�#�%O<�1'L*۳���s�i�N?[��0}��<݁�:��u]�Ɲ�X
("�IB�XCI{�� �}Og���%C�w����q�~��=�
�y`bM�a����N�&��g+����^�@4�@v׿w�ٗ5�<����P�IR����{��k�5�%Kb������xLb��6J]i��z����Ͳ������1��޻�xn�Nu�d:s�xɲu���������27c&����ǀ1 �:�VA�$ןz��]�C�)="C�'{�@`|g�W���=I3(A'���@>�������P��&�2q��}�K��{�H/���@؁ς>�B��f(eD!��OSPΝ�2ϱž0]W�f�ُ�BN����x�`�M�n���h�ӽ|�;q[mo!�R4b�j5l�n{6��i��������g�R21Fv�|oã�a�q=-�V%�r�AC�I�+'z��� ��
o�z?������r�B,��I6�}�����=ꩌ����T�$�a׼[�K��H$ ���T8���g4F[1�1[��b|�Z�̯?��Dae����,r+sZ�rL�0��՘�}i�*P}[O��<�6ט�K�D=w'���|��M�I�����ӭ�³w�V�,QTV,gЛB)����b}�_^�9�?6AN�@�Fi'�+9�C^��<�Wp;�OFd�@�T1�r�M��~�\ַ�>B�A9�b���ܿN�ϫQљ��Y[�l-t�V	�8=ae�.�1^0�� ����2i��,1��r㩴"�`0*`T�2{���5��=�˦ 9��GV7���s��%���o�����}��k�8�f�A�����*$���gL��)ឝ�6m����@�,�A��9*y�'�Ǽ�a����$�P��Z��
4��1�߶��BES[ B�]cs�᝼$���m~�p�����]����Y�"ĚaP=ݘ�� T�ޝ]l�{�� s�1��O��)�$׋�˚���k�|%�6�b6LUhPn"�d���t(�ŭ嫟LkMޗ�.$��	 �$X*�0�'�Rx��|[߫�nq��A}`u݁�&�T���dP�:�G�[b��ҍ�:(Ӄ�[t�Z7$S�,�hO�O#wՐY��u��;�ĝ=�$���$=��S��p��u�Z�5w2}�d7l����I�_u�����'dB}��S�X�����i���2�w ��X��I�n�g� ��e�ӗ�������<��Z1a��߯���~wh֗�#A�D$������m<��O;��V����H�g�8����Y�qg�Q��WL�y;uk�,.^s��h�횚�t�F�X�*����t���h�Аh����T3�e���'��� s�c!�!
���1"u�·�p��Y���
I�)'~XuC�x��M�}h���XC̝͸=�<��ec�<%��Z�ڷڶ���2'�p�aDB�IX��܂9��{�r}4����"�Q],!;�"{����ޓIxH��<͠�_!�A���9a�q��8Y�{l��Ⱦ��:�Z�b�*("*�����c�y��,��2K��]�p����5	���8DM/����(�@0 #�����s�x �l�����j h�7�́N-j��ۇ�	c��ݏ�/����&i7�H{���1�Z���m��{�m-������u�Nf%��<|���LK	�d�y]�Msz�'[��0`�[I�!3�\�u��[�7FCێґ;ɩ{��U�N��Olq�ss/�w6����WԔ�	D (5n���!��幼�_����P�P�"#g�:gi�����c2ͩƠ�rE΢��u�JW� -�c�u��ɌE�xdH�LH+*�鞳AS�n�jw1X�[r�E�*��cE<ǭ�^B���ш���8��C\�k�{0��ݳ �	e��i�m�I[����AHB�� �$����L�ǆ[uX��甍掶�K#��L/{ȸ��<Τf�:�K5��X3o�0�}����܌̯zt}s�|� >��]���k1��_AzX�GGƚ}��juf!P>S��nެB2�!�~�MJ�3A�i�g04�NUN,L�I�C�ƺh����!/�?�o� h�X3�~䦁��M���g��DӦq�|2��/�_'�"܃���Z�if����>��1���u{��6�=���%ظ3��]��H��l=E�#FL�!S��Du��Q�����yjٽ��u6tEC,�x=��r�7�<4� ;{�E��e�u���9��;f�6�*�޶�F#qi��������Җ,�< ��nż�9�ػ���	�,����P�x�������37;;��$�ǟ+��B�j�T�p�a��\�C�"�k�"�N�t݈E<�.6َ���:���:nm��T�����e�h�/A֤�z;�8�'i�۞�M�6�u��n�=�Ϸ9����}���*Kmdې�p�[/cj��	z�����]�W�ܬ%��ݽlކ��9u{EOk��R�\9�u�<����O��s&��Ý�2s���o6��Doag���۩㮃���m�B5+���|;7]�]Xh�mκ�7�:lFz7X�.�����<����6M��#'�b�բ��`vn��3$��&�\m������1���`���U�2J壅��]c��r����ur����|��|VC���V��WU���ٵ��/^}��v��	�4���&��z�smܣ��|1у���'I��p�G����1��0 �c�@���s�\��}��}�gq�s]����9N�}H6�];��@:�e���0����Gw=��D9�`�AF����ǻ���VƖ�n�h��μV�͎ͨ��7�=9M�������M�V�k�cɁݷ0n�"�X��V*�D=\���@vʈ�+��Ǳa�IlsÖGbJ�Sv�NQa�R�����a3�e��'Lq&�1��7m�䰶�UV�2hĹ�.T���UV$TY�(+�:��N�ե�ֳM@%�8��XF[�yY�G��$����3n�(p��3�o�G�Wlăj o{�u-\�m�������7�:�I�7�<�%�?�G�U�0�BvMlؒx�[��ֶ�Ux^��ٹYK[]���i,,��z�e���¸@9�f�j�vwu�����eZ2)�s����<�:����Y�={z�:��EAE���H(�n�����߾�&v�=��,���2;�ċ�Ek����=̥#����n��Y1��f9������}�8��Qɕb���WX��4���GH��ߊ�[�q%�_7k�ߗ�e5��$�e�O~�ڗ�}����������B�oaf�n�&��p��;��Mڈ֊�2(��{���^��;��7���f��d�B�אKP{�x��$p���"k� T�"ʚ�+mU^񄲳�fXz]��L�����W��p��`A�=�����j�����%p��3��n�����$GZ���+�� �ٍ��%k"���l}��\|�EA�9Or��e.�D�DI�Kޱ�w�k��:�LXx�o�=����o�C��(9��i`=c	Q�0w?H�v�"aAQ�{��j���^��>[��a=�(�]�U��XX���ν��˫�w)!�]��6���\S|���[ {�
9��ҝ�C�*�_d��5Ψڽ��g�W��}ݯ��՛���EX�r���p���S���q�9�u����܆݈�8ޥ�]v������kv㫞�Z5m�k������Db"
���6p�kw-��3WZ��6f�?�b�	��ԉxL	�=-� ������o^�2��z���#	}7ï��̒�5�jY�sH\�c��h�}��Aa
:�����8���@:�<k1��O�EJ�$���jG!f��zޗ3~{M���0!��zu��I��mY�u7��w4�I�Xy̱�9�����b��1EX)=	�d�ݬ�����O��	���g��g1�޾������2�f+��:�}l����1�<-�$��c�C;��b��K�%�1�g+7(��`���*|;|��_���gY�X�!�o,�~:��K�oo��}9�A�3����s�^��"��F(�QAE:g�Iۦ��5����@��t]��N�v�������}{�&{�ѯ7�R�*
1��&�c+9�s&{I�l,���y=g��Ƽ���,�ǘx;�m���"�����<P� i�M�ު�Q���n3+��>\g3��k[s��ڨ#"0�VXŝ�+B�4+�8���B� &q\�R��!�BP�icd2���g4��,�N�w�k����0��ws˰d9'Erx�3��J�����>��<%��s�~8g9�u����z�gzܱ#�6��r)�ƛT�O]�0�N�g��9rU")�f���#��ӷ-�W�N��=y�vG�)���p���;���vnM����ţ�M����X���0s�F�Z8�[��V,U�l�f���U#�����$�U32�`�3	?!��f=�|5�d����y��^��;��_]&o�uo@!/��(��۴��΁!���f>��$�׭����`����ib�Hp��g�4���l������i���:Z��o,�bEI��#m������?�v�
VY�Tž��q��tu�r��#"��>�s�Z�� ����Dj��C4�q�,����6�f0���GF��L�,�� 	���C1����֋'�g	�i�v��aȦnu����XOÒ���d�W��
�v:�v� N�K���!:j�� �,|��=2�7&����a��7q.��=H�����M����=��~�'�O���G���ݒ��������|����c�\��O����}7$;�s���a7�9����^�1�%���!�[�Ģ�#p"s*��"�)�g$��2I�=����9u�q!�����x�bZ����Ȩ�"W�J8��4����g����(�ד��������S��?Z3���p5�imڀ�{�<q�~��I|��e���Q+0ͽ�ȹ-�	��t���Lf~��j
��9��
�5�3�4;�HWr�y�xF�H-t�3Ϫ����������}����Pqe�v'�_޳j�͆� �sޠ�;��5پ�^�ش�a�2y򾤰����<L��a�>{�����:R�h[��z�P�Ѥ3�=
��	1
�
B,>Rٙ�(���<.�+|�Ww���U��Cۆ�;;�<D�W,܉��T�w|~��>��|g�y��=��G]�w��o����DDE�k��<�1ҎA�8����e	k�G�ʱ��\!�m�l����)(�KK�ן))]��Q�P�KFX�Ij3��j������S6�m���m ��9��*�w��w�2Aݚ� yqF����~NZ/�>���,ս��[��r��-�P��ja�j�狡=�5�������QDjU����bv.�������(o'1�8��+�m�v��`�X�T�r��5:�{�=��U�9��������D	�M����7�B���x��z��a3���c���H�<.^;���.F��xx]<�dh��s���6�P��e�|��6Z�#:�%5dҐ�ɩn��/^��;���pWZ#'*Q�Лqή�C]rH��z��;���n7]^�����h��t�s��'NhD�**�"<`��(*�4s.f�u	�TZ�Q����%�VG�n��B��͞�r���~����K���}  ���`_�=ݳ|�Rk�� �ٱШz���\���<w-��/b����/.��,pd��l�څ\3`�.bF��  Nb��Vp.�Ԕ��JY�^�u��D_7�0��w��}��[��ֺ�����5�YiW�7��:��8H|g�_]8w(1�k���r�zxֆ3x<���fY� ��r�b��'I��� z���ּ�4��W8�Ԏ*�o�@�E���Y�̖]�����_��+�a��>��@���ԓ����կ�k	�,M�=�;����r�m�ujԃ��)�.�ց:1�r'��c�P$��&(** �n`h ���l�߯���#��P:� >��v����Xk��8]ޚ��۵c�E#e�����(e�t���g�ıp����.Y��]��<��7$nG���R�s�c5C5��x�C.�1<X���������[��nmvE��S�0rd�&��]=y���"�
(�%E�*��˟n����o�)���C��`�
孲���uSXI,ǜ���;����* �M�GCt_h�x���e{�� ��Up.�:ԛ�#���f<-H������D�7K5� 2]�W�y�h, b��T1�C1ʀme�9�v*6R�=-�r��늃obh"]���3�jۓ��m��oM�E��Ϛ8CO;Qիǋ�b��z�9���u�h3=4��`�ۛ��p�k�߮��ȋlջ4��Z����mʊ�D�I%r��\�v�6���a��1�.���p���%�I����=����3�甀/���/�0����8�_�fo� s��<3P �yjD��l�|�k#���cx�@_����(�PP(芝e��1r�<�{��ciY����9��݆�sm�ZPUW

�SPr�B�W'�Ze!V2j�_V�a���~s�<A""5jDDX�C�b��r�u.��@����8�'QL�� \B7,�ф{�/�v;\�J�����d�G @ze9�f�f��,TnևPQ�"�Y�r�jܿ$]��Ր �Q���<������7R�>�Of��3Pr�T�\ޛ���Y����6�6����ڌl��g��"�����`�@���{���x:�9􌇾k\��'^kƨs9���=�^���f����=��`%B��18����7;|����	T��k��OBK��x��oEm��^{o�d���}�ܶWFcRww�� 9sV���O9�)��1n�엗�[^k�y����:��u�8�E�U[JV�mKj��N\�|��ͳ���;����~�bu*�G1��v,*�D�YJ�f����;�^��g<���6��u, ���2[ގ�6���~�1gp۴�����r�x�\�j�gږ�^��G�:��vg�\dƵ���~�ݟߩ�M?ʘ>P=df��*]r{�{$�&.�yɪ�5'e��eR����k�(N��ܸ��^ޚ�7W-�c�L\��v�ዴ���CF7�콈�>>u�yb3Ր�>y��|�����}�;�a~���W����q�==��L�����tL,a���� �U�nҬ�v�<���~�`�/g��"�ط8a^ުY@�8Dŋ,�����_B�"s�7�.��>�oz�� ������{Hx ���S��AI#���m&��K>���b�$j8ыl�q�mi�S���+Ƃ΍q�X���Q���m�qs�q�۳�n��@���B��{d���(X�s�׫v�;)��v3��Z7<��/V�����gn�N\cVwc�|˪�bS����qݶۛ��y鋢��/[�姣6
�v��X'��ޔ��u�u�z��Q֗1n��طe�x=��cژ�u��d��s x��v�
-wm��M��''���V�H�v׍��l��mݤ�6䍹�8y�gAY��<s�n���u�k�B�zz���ۑ�uz��g�#�o<]���B�Tn�`��K)I�,�ٻ�?˼���Ĩ�WE����P�H�������^�5�?f�N$?d�¤8pm���a\�ؐ����2�V��X#pt��%r����=�	"ɑ�ŝDV/t0U�no�YU?5�y��s���꽒{��{N��=�+�D�r�hc��۞�=e1�#3��tw�����0v��wg� &pn���7E��y�<�1�.�96ԦC��{~�I��Y���Cwj�dU���I�T���x�t��N1ٱ���sT���wS����n��|X�D����Z�v[�dG�4i�kC��#�X�F�EZ���%J&�u�㩈��(����ȓ��c�<�c��[��4zx���VCF��'o z�߿[��ˈ��]���``���#��9O'Mk�?��ε�&Rߓ�^�Q�R ZT6�LF�������ߎa$}<j��O'9v�ϧM�=r����	�6��{���/�]L}��KQm�R��}�|[�ʙ���, ^�V��Е��H�	��V�3`Ō�1&<*�Z� �/�>%��}k�%{��7�x��9m�P��pt =��O���F�����Z�u&;L�@��i;��H���v���E��Q�"�2�dD6�V��QU�R���Eej������S}���ya3�9¶�[�}k��O#�,�g�l�+ðEU�p��aId%D��!a׹���0�^E<3�jy�؛|���8���\L�y a	�s#֘��	<� DL3rW7kg^(�lO%��[�,�w��q!��oQB�im�Ym*+W߫���ц��gp��L|�o޾s��Q`���%Љp��T��n�9���ז���
��Sĳ�9̓�86K�� ��U�P��'J�奍�1q��E��xH�>
`�n����OpyE�:��4	����˶�h��<H�b4�*�,�rÅHG~��������ι�M�V�s˴����8�B��	<��1�%:u�y������]v8ڝ�\�k�ݞ(�H�����Vڕ�b+m�V6V6�i4��YW.�� :QZ�W��S������>wsݴ֟��5�4%f@,|y3�\�X���\:	fO>��#uG��z�9b�J�A����5v��B���h�,�s�ew������$Z��:㵯1�STz�r�ϑ�����Hcih��Y��݀���F6--�¬[K
/�}M����C�o3���1��`d�C�<-/�^�����!��N����8*IX��X�jc�+ ��5�[�o0���q��,�4�{��!���f�3���=��x�<�Փ���`[���&Uz�D�L>�I^A$	IBV�ʋb#JR�Qe����f>s���3��c����v7\��&��l�n��w�R����
J�J�a (^����g��sn����e߼���#T�|�Mo'sRo����{�ܒHLMpN"|5�T�:����+�Z陵����m�A@��:�58D@����"��T�jQm�}��zg��[�Ǉ���
ҏGPE% ��K�`�fI���G����'|�c�71L�XRG�2 ˑ�b��7Y���� �V�Ǚ�4��f��~�pȳ9��B�(�QU�5�Hmg�Wl�UM#UnlKr�#F��;�x�����ɤRq� ܯnv���M����0�8-m��;�]9�t��[l�m��狭�k2�N[��`P����)FG��fR�-��jk|֭�� �h��Pm��C�}���	���K�M4t���m�J��D�\F�G���b����f�f�!���s|V���X-~q�v�.�|҃a`@��/d�Sʌ@�? ��O�r~�-��vwy��u���f���ϧ-0�lO[9E3�cY�15QGi�6��Z^D���bV�kU�X����|������wDi�+���F���.�l��#q3��Mk�桛-~�H��R��j��F���A�E'�ZqIGpv���mut���L��2�'�<���@�/y��I��Xt�kA�=��&��9����7J��q���7ٲDV{[E�G�e�a_���jx.�c�'!ڋ=�_8�W���B�K����{H�� �|�n+��I�۷/�W{�����2)��-h�WS��^���^����=��������S�@8�~�_`�²�sϢ��6DC���tc����ܝ>���˺���{}U�v[��9_��muVZ.Ҋ�1�S���ӷv�����l������l^�N/ە{�p�w{!�yN��S��A�wQ��"Y���?f���3u�*A��Y�K]��ίd�����'�u�������J诋�ɓݓ���Z��n�rƮ��c�էG9]���������*8l���fY����=���!&^t���՜��k��׸�k+~ʺ۞�ю��p<wg�T=�Ѹ	�#!IQN��&�g���G��x������@'��w�|y�M9=��߼����I�_K�Q��6ֲ��-��Z�[o]w���2�6�p��$�*=��uy��K;�[�]�/�|��YhH����HYK)\k܌�{�b��^z�i�o��[1'x2�alx;�䋕^������,�`�<CBY�L��n��mz&!�v{�sεފ���ow�9EYPmRU�B�(ԭJ,�^miQ�ruc;��^z�:����� ���c�	��Y%^x�y�������6Ұ�E�>N�3��w�a��w�t�_����S��Հ���!��"���ݹ����"a
8�DsŽ�������w$�
���� M�2VӍ�<箩�x/��[rvsG\�1����z�������7m��>js���}�i�-�N����V"���F�(�%A��DV��ޓk�ժ�Z8��R��H.�Z���@�]�{	fQ߂�G�T��g�ڃ�9�ƥ�����=�0�A�k�s+H�P��|��Nx�Әk۸�租R��J*�1-A�u�u;�cg6����h��,n��Ɔ������8�W���R�y�sݏ�Xs��iPl*
�KA`��iUE-*(���-�ץXDW���3T�g��čs[�(s1��s4���/�_�2I��f'���R�ϧ�"*�&I)d :A�p�d�3�n�w$�Ӊ�I=~4$i@�)�~N�Gr��f7��]�u1����Ly����{U��AB��R�h�eJ-�RإF�;���n��� �h#Lv�Ӌ����gN}J��p�}5��?.�m5���;G$��+����־%oڞ&��Ƭe�cy^���NfI.�y��&�܃����n��17L-�2�*.�l�\!ͣ�7�i��� Y�kF�-EmK[B�4�����	<	7�Hij<2��f�K!�H�X�����m�KU7����4߃�n�*�fG�x3����FC���E�
�v�fp��,dk�X�g1�X
�c��b�s�;I�Ι06�\͸wyW2�e^�s���P/��d�]�^�Ok�h��G��W�a�ֱ^8�V<�c�����8`k��uc����"%-P .*��J��Yo��jEUlux�3/��a�eI�V���o����6���8�H��`�6 �m���ґ��I=Y�M��O���{����Is���k�� J
y��L��OFxC{�1���C����zZ�:�V�:).�s$���og��Fcg��)����y�#B�i����_�^�z��mM�خz�m��YX�Rߵ��w���LD<��c�3*�25l�fw�N�g<;���6'3�s��}��<���Kzz�f״���^r��&��
Yde����y{o�gv�>aY����i�F�g�Ի�� L8vP�y��]9���Ybj������e���1m��l��Ɗ�Ȣ�U�YF0��z��e���C����≂����XXЍ̞�mn�,�(ׂኩ�23��`Bщ���b��}kˌ�,Wl�|�%�g��BTQ0U�H��pg0l$^Z�~�l�bGI3�TA���¦Y��q��-�7z0��8b\���{�k��=g���}v�z�E�Z"��
%��X5(��[Ϩ���$��־%�Q�8��q��}󞢁mV�l����(ѽ�8���!�eN�˻��<��p��EGOa,�߽n���/h덠_O�iw��Qt�V��ky$�zَ�,L,�[��+���\�Eš0��8U������fʨ^�c��g(��}g�p�����'�����$������sq��6&���ޏb��<�8߁����QV�N����G/I�.O f撄��=���?hC;x\=����?<�w����^�쿢�̹�lõ|���3�,YIY�3���
_h��G{;�OХ���N�0ŗi'.�V&x�����V~���Y�3����=�͙�"�O�\Vmy}�=����7�s�R��TwrdZ/����򴙗0)�v���z�\�C<�۷:X!�h{��8�j�#���,��c�U5������u�z���wc��&��	�g�c���u�vI{b�{c��3�@��l'n۷)��\�p�����cq��`{�+٬*#��GZ+���x��wZ-Y�X��ݺ���s���@�j�o!#�[	��T��S�z܆�Y��xs�����K�۞Ne�l<�tm/�űc���v�uݫ��å�&ٞ�6;;���v��#*ay7u��<c[[��퐲������Ƹ:x(ض]N����M"�Aз��7G2�Y�D��ćj'[��Cu~��܇Y�����7Ţ|tsh�z�gznQ�K�fL���&��b��8�@SoEU�a�,�ʲ�� �Y��
�g3۸��ם��G���~6�
�_�k�Ax��W<Wݛ;Nygxx�����;v`��Y���=�O9��nL	w>�k;�A���7�t���r�Oz�w=��f��}����W�{��{��������N��%Q���m��J7f�Eb�� ��]�p���^�.�-��3��;yx�v6�x6�3���Q�̈́9�5�=��Ϊ]!5�����뭺������+X�QF�DKUV
���`�-�J��4��ֵ]B����DW(�,Gxֳ>��l��2�(������lǊ.�2�z�w[�X�Bq9�Ō${��n;��r�4�����dt�6�@ݭ�%�`�-@�����u�n�����J7,x;��k�1Ѣa<��M)�LԔ7*k����O�lX�j�j�
5�Qmib ��д(����*B��k}�}�	_�3��L��(A�^;���3�[ b�����%ܟu]� �6�1�h�d�8�vix�!�	m����Ȋ$���moϘ���[�Dѭ?9�3c���.�0g��P�1��X�5��[���>���wOG��CiR�����}��DVU�d.Z�1XT�������\l�ܳ!,$"��	!���2� w4��Rj�@�����$��P�/�]g	�V�*����&��p�8��3f0h����W�B�����Y��w�J��Ģ��ˋH�=r�����z�bx�����n��,j�6�`�TJ��=����o��/Z,(�ZTb")V��/�q��̵*�Q�.R�"ˍƗ+u����k�~k�ͯ����if�I��J�c��n�2,��&i���`��^���e�L��ޭ��4 /fe�x�O
�'7k��T83�{�����^4�pg�"�6��]�.�{5�����~�is��m����^�>&���A[�p�
ۋ���vl�\��R��v���x���n95kg�u�X�M2x����eS�J�X��b���+Ko�ڦզ8�F�FV�L�J�Sj�^mȜ4kd�#`����:ۃ�c��^r��3�w��Ʃ�J7��C���y�k�;9�9�ܷ�4��`�D-�>��g��(�p������i)���{Q�m-��$$"��Vz�yq��+7���}�N�c��D-�|E����a��/�]������:DL͙j�R�R$q0$*bf
��ԩl�TQ�[k(H�Q�-$;,����S�x�&l7b�]�ji�d��.�����!���:.�7Әު�_8K��8��)]u��Q���"���k���&���K�����O�@#x+�ܢT�s�FՓ14������H�wy�Xw2"�0:�(�`���TLDr�ԫJ�Z�Z�[Î$�y�<��o4Js v��*GT�K�m{S�����o�
0j@J��LF��(����5=�$��j%��G[��c��2�7���X��.Mo'g!���a�(U�QcR��5
*��բ����9MlI2A��O"�2��h�e���̘�'��]��#|"�>) m��
g"!h� !m
��%�^f�}�&G�o��o`0��� 7Y�䝜�Zl������`�~Ъ]�@]�ݲ�#���~�"F��q�Nvy��kqb��scX��af����)�:LՒ�7& {I�ۑ��ۂ���t���s���d�`�֎���4�p=���ۓ)�v�y��Ͽ?`�mǳ)iiR������[Ym�Tiݍ����}���V.��ئp]߄�d(�����5�+��o-�gG%X�&��C׼��1P}�/�=�is���c���, ��#ٸW�o�WZ��h�n�1���D`C�y�B��y�Q�U�Fr��=9�Y��_gZK�15��*��'	$e*��J�-"+Z��"*�]ڲT��ren��7@W�G4,x�J+��0�>�b��;�y��ϋޝ��1�s�Y�����J@#� ��A;���h�^�ݖ�s�ƾ�H"�v��"�dߏ@hs��ɹ4Azq�&Hz��̋���vp8��̙��24\�}��2FʋZr���$�[Z�k��/�kv���<"��.ǀ�����Y�UH#ыȽ|�q�]�L��n�E1����Ѿ�U@g����k�'�i������M�w����r-�?cÔ69����uqwџ�%�F�N�w��8|���_׶��ی�[��6�ZӸ�`��b�t
t0���x�S�}�l���,{)t��֍�?Rz�=�8�*�4��(ȕ��VEP�k��Ī���ݤ���`��P�LB�O�rf�����7�w��W�z6���%���u݌;�*n�5�y=���r�2*��n�N�~���P\���=�ꏽE�Ӳ�G�%x'#��G���x ���'S(O[����ߞ����)�,��+��}���v���������/_e�Č���>���%�fC�	�X��+(�^+5��R}�5���x�:a�#��}w@ѿUZR�m*�5����/r����^=����)�<���Η7&��ܨ@5P�:iB���M�鎃��w��5�?���'�[=kP�n�2ڔ;����sx����fܽh$~��ϲ6a63�~��4e�"VZ�U��Z�e����͟)��w��ϯD��Yޙ	(0���X��-e9�m-���riu��xC�U�9UCE �i��ax�{��s;�%�������{�4�H�M��Oѩ�س<���p��LG1+�;Wj���;U<�7�����`u:}����K�H�M�;�C�g�nG���s�SWX.R���|�(�"�-��Ns{y�Er����M�W_��1���_x�wso�f���wM�\��v�/a7��h�:�2o�5�˨ڏ�o��J�^]!h�Uo�>5{�v��z(b��G6x|�}�Az������Ȋ$Z	y"	D�" ���W6 Qє��eC�K��{�3��rr;�J_R�r�G�v�OjB������@v�A��X�N�w*<�?�:X�g������w�i*6Ӛ��{`�s#M�&��aY���q��ך�kiZ1�b)J)kFW����������Z��vky�up������]�FF���p���V�Ud��]_,/�Xk��@#Z~s�)��o�K>�@]h6�l��<q�f��=��2���n�f�5c�t�Y�s4�N>���0���R�5-����~�)��k7����3i��I{8�5���m�TJ±4��݄��s��Q��S�x��5K���;E�#�<���h#�����]0<j�=C�`�;��{%���J��C��.*#�9�X����en�^�%�I���(SNN]'[We9^��S��L����b�lv�U��ۭÐl��u��n&GG��[J�YZ(�����O*�qƦ	<`n�7C���h�B82�\uг��������i(+�m���u���������K;�Y���m�
��#�DMdds�������^�T�c�Z�,��������v���KP��r����oz���\�Z�m[(V�>)5�
"�g��N�E�`ܨ���N�
���u��և��M�w��"�YIx[r/=�\a
9Z����L;�s=�*���Vy�GR����������`�dL��� ��M
c����f�F��p�*_�VH��r�-�o�*'�P�h�+i+O��F���p����!.A�x�]�Z������Z�,�T�\����K0yxU����nKq�k	<i�pjl
=#g��2��=�.��H�>D��^���l]&�w74f��w����ҭ� p�����/�� '��>�� �
�Q[bZ���*#{ߙ�m�q_���wp����		"�E(�@��nT�>�;�Y�0�9�ݽ�.����O	��u�pd���ݺf����� W4���6Z;[�w�>�[ɭt6Cv���s�k�.Vv�����
͛�T��{��݆^��{L��m�܂r�V����n%=���Yh�j�n=�PM|p����j������#��'x�P�<��� ���b����{�zOz��_ocu����q��˃s`��+AY��e٨Bە-*I(Y*K�nj�U�9mm��9�g:7��g,`={Rժ�����|�9 ��Zß����A��^�a<흯��d-w��~�"D�]��zh�Y >`���{�����5~� �Ɵ��]��9�l2��o=����;�G�'T�ᕑx�xܰ<��*z-����d�#�xu���ۅ�[+�;�+���5�0��U���gv�<�mƹ�^�!�^��^Σ�M�vK��疸�ȝ6,�p/X�[�6�KX�6��v7��w��E2����1���z����1q7"5Oh
�.O�C�;n˵�W9x���P�4:*����Pj)�5
�:��t.2��M���{�� ћ�����nH�v�v���o���۫��MΧt�凲kw]N�9`;j+z��xܹ"�ֳ¼9	�:
a�)�=t���m��]����V���z�/i�W�?��'�~/��˻�Z�t�[���<�����MǗ�jۇ\�J����i]T��3�Oy?�*��宎O{z4�P���8-x��VX&��s%x�Vd)�x�^������z)�w���1t�Dg#���Q���|�n7�ҭ�A)Ƞ@z�/-�wQ�G�����幃��S�{��M>�v�ZOg������M����}w�f%��f����}�xZ�y�c�z��}I��vS�a�n2�k*Mח��c�Sp�t�L�\�;�M�G]�3�V�t������-Vfٗ�e�k�Ԙ��{���Z֭,j����`�YR=i�0�V�mJ8�AUJ����������o��8<-����n'���RE����]f��v�T��\7h�7 ���M���W33S����E���X�YTELw�x��]��g\�X���A�!��OX���y5����=���t�Q�kF�6�J��ڧǞu�@\����n��z:�s\��^��/��𮀹�f�	����o|^ݶ�Gh�-�PpDtC$�ü��>��1Er%P��s�1K�[���2��ϻ¾��Y�CgEOR�+�٦�*,��	����H^%��X�����k-���M�G�n�>�9�x�3Mw+w����{�B�Sd����zZ�:��k��抿����y�q�D�2x�D.�dH�@7�ɝ_�3���b��uJ5�m��N&��m�7��s-�C�Hz��QRҖ�A��}����o��7��ωża�N/K~�bt��¢\R[IkP�=�j�KbmyysKpxڿ�@S?��g��Ǐp[	�ܰ�^,;����1���`��� #9�-�s��k����j�W��kokX����;�5��*�	E�A`�nb\#�`MK�v�dG[�/l��t�7#[�Î;s�1���i�;j:^�ݹ�ه���D�G��
�iVڻ3X�F���aG!+E
{ݙ��� �'�K���>�Uq��<�T8;�bW��m�ބ� �Ds�ȗ����/>�����l�&
�Y\��+�+�{��B��@UH�����~��Y�Y2�z���e[\(�YC<��E���x�(��ʫ�r���欄o��;��No�s���H�2���+�4y��u,�>��@��ҹ�:I��{GQHȪ(�
8Q�E����l�W���+�S��<8e�N�e�R���7��Z�X�P��ͭ�Ӫ�B�j�jإ�U�/����::ַ�x�R��W�7��^<+�혞����7O7.Yk�e��0z^���H���*�h���� �z�k��9�ڞ�T����2�M�:�y��Ds~�B�p�wI�\�;f���������DPAh�k��n�|v�}��Nicz����LA` )#���Y"�]��G��fw������_����fl�v�O�ي)3�����{�_�ρ^ގJ�;���C�O?T���:�ܞ~�pY��3��>L�w�Q�T��IJ��+E��ؤ��:����Z[ut��q�\�.8�[�r�ct��p�d�v��yƼ�]n����v�+TF��"��*R��~?�\�=N;P�Ft��������8_aN��io����*�6b���~.���Xވ����~�Y;,YM��EAc�0r����uvp��2���g��;SMyLÐl6�l�D�ȑ���_"RA���$�Z�
*TR҉�}�;���sϳ]O5ڝI��������N��gɿS�nxg�U�0J6����H��;m�K���xx, a�y��^�uQ�ȞF�}g��!������a��_�mGs�bĚ�o�hu��f�h7%��懞�=+��7N?��_h	e��W/�b��h�{\��������,�8I�lWGvF��{7%y��J���s��.�n��'��U�j�(��a���.��p�Ž���qOM��O|8�Jؽq�j��~W۸��2T��
��
/�x�r���c� �1M��=�;�&�����Z���j����n��ʟ���������ᓁn]�TZc,�3�.�j3Vyκ��!5��j�W�]5���wg}�J��w"b�Qv�Tg�q{��{�}�=����[��@RoOf���������}����>*��gFy�aq�&�(�����̏o\�O/��P���巐g�_y����+v�8$����z�G7.�����}��*�t����w*�w?wn��6�{#t��=�;d��מ8�ց�݌}ݜ9�t?S|�z���X;4y_7f��;@��7�5n���p^ه���'�fӝl��C�{���;��g<�~o�����J�J6�]{2���a'����K;�y;}+���0�|��蜒�*�(Ȉ:J��B���fp�I>=�fO;9h��o�uy���!;��f������.���x�*���A��g�{I�5Sl�2����1u2�H�H!� z|zx{�������2�O}�d��%tl�B-�_ve��6'�<�ǯ���n��>�5���������D�ۭ��1S�C�4u.����Zׁmv�;�3`��0ӳ5�L�~�H��z��UV�B�F�ʤsq�|v�ckN�ós�ci9s�G[����C�[upe�8��38p�֥��Ʃ���AA�"&�n�ݺ�'�[t�ec���vo��%6�Qt�ե�`��g����
8�e�h
u3�y��_��L!ܫލh�>`K� ��>�X�}�w��E�WQJ+�d����z��T���ə㷜l�;c��&O,g��v�0�7�ޯ�3x(�骭hϯ�=�:�&�;&(���+Do�P�.��wQ�垤ܦ���y*kA��
BV	�"��K���F�q�<�w+��g�t� �(n�k$�^L�xT�����}c5j�fRgڅA��1ٝ��$B � aiW8�·�Z<}ʇ;���U)�ǑU��Tp�E	l�2���/{�y�gA+��x�~4s�C��z1��, ����Q��W��9�Ι	�K�؃u�D��-	�e�T?��5����0v�DJ�+KQ��-�m��o��$�>z������V%$���B�)J�tat�l]��s���+�P��k�3&g�)�z����y�����N=XѢ��A�q����=]s��G�̴�݅��1A����##S2YwS����!��P�;\[
c�8��É2S�uq��j�����	���0�	���[��n--��\p�bڻ{�`�%�PUy�m�p�.��ҔU�	P hT�7����aSqyysb�F�τ��6���"�4+�ӎ�Ms`x���u��лL�4�7Vz��P8?�߶�K�X���T��d��E;��ŀ�P$p湣��+|�fTG��?��:D�{ã��8����0`	�(ե���|ߤ���[�jf�<�����N}�ˮ��sS�s�L6�We��DK{�;�>GA�8����L��R�|�{Ė��k�~��s	�ZClӬ���7SB�=�g`W-�l�A�*�\E<Ķ�a[�90O� ��*LEm3�T�ݲ�~[x�˄ON�<��ě>�X\y�Q��W�L��K`�B ��[��s/8����rG����Bq�Et�4D�)ucܽ��T��L�n�&��25k�ow��ھ��Z�A���S�nd/Q@����@�]�r���Cib�c�;�;� ���L���Q2���5���JG3��9mB�qd�ƒ���㰮z	]$�{ӰuǄֹ�nb����W-���>���c3oF�m��e�"p�}����?F���;~���M�l	%���t���@+$L���1V�8h���4͊[5�l��-�$�mIfDڌ� lJ�U�Q�j�mU���ʎX��f��JleN6�\hGQ���.#b�|��۫�MI�"mJؕ��̀:t�ܢUt�T�MEƣ��\$9���m�sk��Ķ�m��L�ቴ�NM.0��8���cIl�V�rj���[P�m\��&�Z�lmJlڪ�N3h��$����n*�����#N�\��ۯ��ٽة�HY�L}<8�~�3����vu{]�~�_�������?����'�r��g�q<Yם�������������=G!��n����>gONӅ��=gy���N��x<H"{O�X�<}g�����'�s�s�PD� ���cp���}&>׽���]�Y�����y{�y�,���o�^O�@����^ߋN��g��_&��?'ms���Ε�}�Ç����e8�qӧW_N�}��t3��'�q�q�������'SD�M10�2�1�d���ȍ����kR�F�Md̪�S04i2ԙa2�5jMV��FS+Je�0`a�a�h�4h��U��1�jԚ1L�L��S�jM&�SE��4c#[�5�Z����45L`�S�KK����cL��S1�Ʀ2kC1��V11�Ɔ5X��V25����F5�Ɔ5�cI��Ldc#��Ɠ��Ʀ4kQ��i1���Ɩ5Lj1�ƋZ,h��ƥ�V4��c%�,dcX����bc4��1�c��1��h1�cV4Lj�j�j�h1�cA�K���V11���k#X���ii��XɌ�j5��X����V0�dƫ5���,j�e1��F24ōV���ƣ��2���,bc%�,di�cI�11��+4ұ��4X�ƕ��&���1��+M5j�`1�ʍj,d��X�X�c*Ʃ�+�a�Z��,ccV��M5Zֵ�c,i������kYc1�c��1��mKj���V�ò�q��X��V��VT�I���Q|��p4��ϯ@�L��7�{��9_e'g�a���|=�����g��ud��ίeƻ��������A�v�s�'�����:��z1��D������u�/������/��f9�i��?�r��>�r/>�i>]�^��t����4������;������a�P"z�1U����z㹿Y�=��߫w|ӥjt�=��Iչ>JO��}�j�/��a�o#��}A�|O+����#�����N�������;K,���.�����o.Wo+�pU��]F�+��lss8:��e�s�Dܰ�:��~I7��΁�9�W��^����~c�;���|<���3ʹ����t��/i��O}����Ok��|��v��"n�|��?q�>�t����w�z��������ҹ�6�w#���n'&�ܝ�v���u5���z��˳����x9�r��ޯ�����W��<np���,��./����z�y']C���f����C����tS���ѥ���p>#κ�="�ӝ�����vD��ns����=����xc��������uˇ���r�9��{�?p��)�����