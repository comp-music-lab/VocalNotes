BZh91AY&SY"Bxp�߀py����������a�?` P  P(            �          (  @  �E
*
**U@�$�Q$��R��QU"B�JR���H�T��RT�E%*TU"��A!B���ATR�D�(  �Q%    �"� 
  ( 
	 �T��
�7z�UD�BTRT���ȒB�(T�&܅��9 i�\�B�l`���t�PV� ͇	R�RP
PB >��վ�A}>��X:g��D�J�\�>�WH:Þ�.���ݡ�t�OM��S0�/Y�[��z�N�W����gZ�%RB*�=H(�����@�  hs�#���r�����A���<m;��ZT��UI|M�R���w�;҇͟M��=�>mJ����}o�hc�E&���M���=1i}�Q*���  x�����|{��qECrT<-x���/]i�H\.�owR�<��iꡜ���Ҵ<\�S����t/=�G��=�t�U
�H%��	T*�HTB��R�@��>3|��u]ͪ��}���� �� C�6pg����vy�{��0A�\s� �"�T��(^C�'� �R���9�@;�����@⤼���w0>��4�`��TJ���(�$*@
!.@P;��xA�;��vvw`i��@���ÐN�ӎ@�����{!HT�JH@	W@������� 5HK �@��t7`����^[�2A���a��݀��"�[��P�)D*���� P��^����1W0�0 �zP�g �9�=�;�ɈM�A^��@݁�R��D���U����8��i�8���{���9 ��v8 �����=��|           �@  T�2R�$`	�� �	�S�a%)U4i��421�`&� i��4�j�FR�mLFF&@ d 6J�&J�ڍ�2d2 `�A�	OԩMTр0     %S5U!�4�zCF��
{TcH�S����'�~
������X����ҿq�}�u15�w���QPAz��3�*� �@QQ�DDAb������F?��������~$`�R��D��|��� P[b' ?�a� �/&"��~������(( ��d���,�c� ~z�<?�!���?�R����?�_��I��YND'0�@��U,}��q�ռ� ��݁|zCu�Τ�'o>9�O;�d�vq�Gw�m�룯c�qU��R��Ny�f	[�ڥ�@�Fu�jU��9\��5Ty�3x�z\Wo&�l���I�v�y� w�:�k�(6qpeEϜ�Y[�m�ܷ�����G�s���I ��j�ݧ���V.o۷s�s\�r{z\-�rް��:u���Z�Gh���x-|L���X�|�s\�k+]��@����l��B�;�3��gt�yw7�`
��>qg��ݯ�������U�s��z���3zkլ�G����n�G�w��@X�#��vn�k��X�4����EZN7F�,r�b
�(0��nwb���ÏE��hU���+�Rx�Cg
�"g	���Cǫ�w�w�e>=P}�γG,6K9�N���.��p���Z7o	�OŃ"Z��c��1����m�b��9��:N
W�nKP��u�X�T<�����/c(w�/[�+��� Q^����vْ��ߟ]PS3��j��rsn��ۏS�op��6�QW�@O7F1f���v��'������;�$�wm�:nRW^�Wh��p[8]k.-�V=��c��K��tq¡0�櫡^��NۋM�1,8n��P�|�(ޒnj��')oD���%!��^��G$d�W[�\�%���麳��W���9�9-'t݄v�k�V�ZY���2�������C�:Xњ��� L��oz����F0WN��Ϯ���6�G���MV�ۘhR��ӰQ-xct-l��}Fl�r-����Ռ(L��d�"[8�/8�^wvmK$}�C�Y�5��n�<��&`�o5d�]>|�H����Zi��t���*F<���؃ WF7���g7�x��ʡ�����	{JI�{5|��БW��3�s*���gl`�j]�E�Zv�k���̢��đ�P��l��^`ńa����h:;��\��79���{)����lwx�_�`����M���b��v�GHf,�P�qmjc�@"n��������0�6�l��:�>`�p=z]9)��������}p��2
;Ӛ�o�tj�̧"(^őќ����U�	�{' wX��7����ge�����bg8�+��o6^���!x�w{1�Q |��,�]t�}�s��������NH�|�H�R��N��,wJC���p��7�0�1��n�0S�1h"�Ӧ�d��Zs������ٚ�8s�rS�ebǭ3��Q�v�nTp�Î�aa�Bdc�gm0�&<���J��">]�9X�{a�0�� 	���T��K������໴k�X5���A0�rei&�j��r� 9WN`i�#�Ο�N^�8��oB֪�`��;�+vQ@e� �f���DP�8�H�.�H�[�ֳ�R��,y&�VP�Dѝ��^�u�s�����}�,Y�T�S=q��q0r�ی���7���জ]��e��qєnq�D��7�E�9�oL��٦w
 �!٣�T�i��u����U�����2�'erF��l�׷��3.����Du��-Ǩ�K",IǛ�������uc�o�:�ڷ`�p�q�͝f���Hg�Ǌ;�rQʾZMC�P;���4�X�M�R	sw�]��2M���M.�;q4���ۺVC�������ZΪ�u:��ծǝ��Y7��3B�Wë�/px�����Z�t����5����x�#�_�6���}��7T�/����˛F���Xtv�I��03����2=/��!��{#�����{ٌw1�쌫œ�o���it���Æt�WH�M�nu�����!��0��s�,氾��-��"�)1��ׇ��HZ!f4����,Y8rf��n�=~�{9{B<��T�w�G��ggn�r��є��ם��IHrE'\��ͪ&tK{4�������q�ٷ����@clk����c����D��� [�p�L��ZZ��7�w���,�؟����si��h ����`�[���Mת�.�o5��j����!P�i�@����7���K�«؍���V�,6w,�ґ9�({�;qn�Qдo\D�� l�Q�&k�4�m{s�g=j��kЊ�/���Y�ư7�����8,���N�9wV/�hrm^�[7�o7I�tcmkQ�.oɑ�8�7��,sHȖ.���cΜIڻF�-�WU;�sEx�]��˛����.�;l�нY��ø0��ᕌݛ6�k^kϽ��ٷ:��o�k��'�����H�JV^�m&�V��ڤ�	<'q�j��E4i跏p��nۼ^�u� 9wc+~����K��kq�CB� �`�8-:+�pj��[�j'����ܦ�4���g�i��<���:��/[�Զ�s��&���	���ˁ����r��z�Br �<�Ԫ��ų)u��vLNK��V2��Kv�FI'>�ռ��$h�n�gK����� �����ӄ�S;��{�vv�c�ɡV��!���?)�.j�#an�(�w/�o�)��oɺ3�<'��갂z���M
[�������]L��)�а."5�>�4ن�R�&��ȍ��������5���q/�Bp셧���hX&^I��a7N&a+km�R=�8���W�j�y܁&p{��!��U��0q��r��;�Ѭ-�=<*��v(~�ݶ�s::��ce6-#e5�k�;p��ޒgw����1�õ���{@5���sL`>٫h�vjKR���ה͵�H����Whv��8Zz'N��<\��s�TCxض�{�m -��ǑSy��v��F��Kl9��s�#ɻ�g�'�`�ֽsy'��ŵ���:I�@�r��w6�zY�$�&Ř��Rzz�:�!oË�;�� �'���uq�Rٱa�!��i���l�f�����9��0j�4�wv$ˋ��[���/7^��%���,c��4���ڰW�W$��cYl�oZ�
Un�\ۤak��3�*>�t몂N�Cs�����hY�l���X�T���m*̼���d�
-D��oa�Lސ	/��aô�D�^�L�-vE�wpޮ�����{��]tm�rB�E�ğEԌ�j�0�k�@�Uʘ��
=�2��J;�{�;�����ml� �l���ݐ��m.����j���#Ӕ���T�u��/Pk��C���F*�!@���T��܄�픽��Al/j�q��xv����'S��F��vͭ�Å�D�r�޸���������I��G���J���3a(����p���!�2��L��=�N=�d�'5���;N�[��w���&��k�$��W�F��L�ۛ{������~=.YR;��7�&��t}����Mhv=�ʡ���+��$�H�<Cw.-�7o6$e�D�no�ĺ��6���EYjc��=�y^�ID���̻�.�$�e����Hܵ���= �U�a"P$�n���I`X�w6��!��!�w���V�$��݊2�G	�9���L�x��ŧ�X�]���Xnn5l ���t�X������c]dj=�����CI���g��9�ۮ��n
gh'y.��N��hKi'(�4ݎ�2�ۋ���Ӈ���lav��!a�Jr�g�O9��z�Y�:"5�:Vu���\h[��;�k4�\�ap��yu���{wAޗRm�іn܇NBs{���p5���1o�H���\���Ɩ�N-�plv]�U�%�!ũR���r%�����{se l�n6�ݪ1�mI��7�B���ˇy&��a��n�I�w5c��ut���k���5�8�C�p�}��Ý��;�u�O\�ZR�ptc~Z�Z���He���Ɓ��Ŗ�u�k�+���D�Aҩ���͈�>��nZ��5��̼1���'{�¯�:�q�q��DD|��׋�N�����2,rG@�HDI�9�Ӌ�Xi�-�����ȃ'��r��n,�����K���V)��'����fv>�����^V�7��X^�y�fM͕j�"�W�N����t��C��r=BY�[ݦ�'r;�I�&�wVl4<'"��	8C��Y����˚�����#��ŭ�ݝ��ˮ���bj2��.�Rx�*$n�*3Lx������GpUK%�0��5.�7W�wr�6�,\*;݉܄�ȻwQVl��}z�V58��WM�;N�
a�5�4��wP8S�p��d��R��Ll��=�^��;4gM1U��]-��A�7��֙��&ps��N�Zk<$���w�Ɔ�jH��K�A�Ϫ��e�1t����yӢ��½�7wudM�4�&(von� ����s��KѺ1�y���C�\]���Bn�EM��8E�xH3�s@����F��B+Lv�-�r3��D$�L�]�uI���N�yLs�:���t�Q-�gQ�ؚ�V2�B�(nͻ=�K���1��ۏyb,����r�{v��1�,������θ�+ �x\��+�fu�%��kzwK�¢�q�q�V�݇:Y%h;�nv@K��4��Aw����p��g19�ws*��Z���kc�a������0�-�K����B�wכ"����G]��4q!��>�0v��g(0+�u=�n���4`ɯzk��<HV �(��u��r;����U�@o�����b:k�iʡ:z�B�x��n� ����/!��;\/V-v,t�U��N���)���g}WCP]Өgf=J�̚�74g�qׂצ�Zʭ�r�%gY�Y�=�~
���<[���?�QU��cGL.I�Շ�s�ƪF�OSчװ��*<�X�7�2pћ�w4��9(5-��2��<�+��9�5ܮ�u�Ӛ�]�D�@W�N�Gi\��~�o1����L]�7�:�*Ǐ幺j娝�Y�����px��~�F��sk�u�.�ܸ/���ޒ�Ҷ�7�9d�/��J���v�ON])�n�������P�J�J�F%J�2&�b�Z٭��B�����<ځ��N�L�t���S���v�'\���q����G�-�@޺�b�5v��I���(�Ub�;���{Wr����Y�����`�4���*$����N孙Y�e77 �2!��L��!���a8J��Ai�����^i�1�o�t͎�Ժf�6GGs�e��o|1�g���+��c��ۜ:c�;�-��F�6���I�
:{:3�7wY	�qO:V�.U�I�J��|4.��gt%��,��R�Xr�H�������քo��Hc0�.�������.�$���i�OZQ�ċ�)�����Qt�C�+Z/��ܱ,�YNKWH��d��(���3McE,˺���|�sSX��ZwTxvc�<��򭷴���ǵ\驭E\��/Tg9ˤeǻw�l��2t�3�aqS6��|�&r���89�Z�Yd�4�r�x�P���P�ꥍ�[���7�`5�͆�U0B�̂7pF�!왧F��jrgg]ы�Da,L����'�l��<;�M��ڂj�S���Dn�S���˹ �aީ��[��_��L�.	��3%�5�J�0ףok�dt���N�J��j1�y0Y��F�@K�N��;��/���A��Qr��0J8�
vk���7�a��p���,l�N�����lwY�>�*G5�w�]{a��-�u.1"���ǂ�[[�n�R�]]�ɖWmԕ�vh�8N���Lw����6��J ܀B&�K&�ti�oBE2�X֥��^W(#E�B:{#�G�c6wL�o3��B�]I���)�)���|��%ޗt5�w:pNy��7W^%�6��\1U3�	�w{tG�Gd���6�25��OP�
<��GwS7F��]�)qq��d������@�\�n��7f���x��<��_R&�c�Dl�ć:���k+F�Ƣ��a,k�;�c79�nFu+s��Z��@�o�ō�.��^���ln�eO�p�6�ܖYc�`���R9����tP*V�gI&����^%z#-��z��A�Y��8cHͤu�h�6�D<��Z�Z�f�sf�� Yx���G*k!�f�ư��uI��Th�n�����M�N��!�p���qn�S4������F�11�~�K����0�ߨ����?/��_\1�����~��'�B}���g)�æ
qN�.�6���n�Xn6�7(���=1�XIv�Ӊj3h���J������ �C��bCRm0�Hh#�B3��F�g����dQ�֖�Q��f��kJ���	�È-i�&h�Xg+T؎v�V�jݵo���!
���v]�T��D1��t�4�)�iV�\[c nXɘ��E^��cJ�̃�-�RQ��Y��LE���Z(��F��1��Ժ,��Tea�X��]PB�(�s)Xe�h�4l-�x�:�,X둹DɅ�EY�*�!���&�=�3H���U6�nj#l��Q e����78��aVD�J[(�<J�܍[-D6���9�,#f-��)��jE1�&��1���+���M���K�SK�ˋv�-%��ƦsUtD�6��v�^�D4�p�7l�.�Z��ie�h���9:��@����Z���j9V�&�%31J�lҪDqu�)����W;@�!�wm-�p�f�&��s��[@���ŷv�M�KJ奶��/QA̔�B����#s���#�
R��O|�i1ڻ V��h�m�`%e��\4e�c���Ř�#���l�-l`��v��Y�a"991wRkU�Xl�s�������jJ6d�|��/���j���e����nQ-��4���G`iMv,���*\�rj�"R��QXMV��w��R�l��fn#3tA�ո�بf�c�6��&lk4�ZZ��&��Jb��v��c�@!�*��hA&��YHf`6�e���VY�!� �;p��u�0+�ػ�vItU"��Ōe��1su(��m��L��!�Q����a�̥u�ihQ�굊�5MtƦ���j�z�c�
LbB lWe�#�M�h��\��tWf@�Q��J�-��+a-(�+��,�nұ�)����644��6XP��`��elo]��F�w���6�C�*8��\=`�R��<�m�vFP j��P���YlK	b�ȣxж+u։��i�:k�˒k�l��aFZ�нz��������5����\m��.��� �µ���X�60L�2�g����f�óHRR�i�t�AK��4Z�p��0` ���4��%������F�m��뱌�c2��r��R�yz�.�m���T�ƨ`G9s���,�싱�9�c��	fьҚ�̓a��cx�ܢX�ĺ1f��Ri��1XU��D�Q�I����(F:ݚC78:�-,j��L���<͔�0J]IX$�sE@iiuԶ܈6R.�9�����f�eEħ9%�����Z2��Ɋ��lVhDK��V��c6o9ؘԻ73M
�fҦ@^�c�1�:Z��)5�1�Ku��u�(h5���٦��`�8���¤�����)m�ݰ�L�p�jG��\��M~<���6��L�p#yΚ�Ac���iuQث.�Ǆ���.���]61oi-�*�TMj\��� �鵈�o()N]R�m�fq��i��4�qJle��&� \�J��Z"�%h۫�,��YHL'j@˛a�~:�ŎR.�љ��	se$J&fn�.#IaU����Ta2�0&5" �@�q�+`%���v��԰�G15��a*�W1�f��Z� T:ܚ����m)�ai���S Ue1�*���`5�0X+�ښ�m�Q��U����[)6,#Y���:X�J&y�T�[����c`y5�e��S�8��c���r��l�\6*.VE��R�`�i1p�����0�&P�&׍k�#{a�j�]�c�m�ٰ�d����X�՞��Ĩ��H�"Jݕ����Ŵ�
l��Z&��-���dnԙ�0��iaF�u����f�-�-ni[V4�c�5.c!�b�i��.L��H��4�Ƴ#�m����ZR^�;��XZ���1�9�n��#���9�Z�^��2K��XA6-��3��&l	�fn�B������[�����Fg����FY�bV�Bl�c`8n,a,� �PѶ��`����Vn\La�uP)me)�d���n�u�
�
��f�z��Q�T�i4�f-����&�Z[l��l��l�aJhP��%i��M0�)���h6��UYY�l쑪�M�L�͂F��lu�[M����Bl֒��tM�C�5�t�]<�j+�J�!�k�	w
�q��(kY���T�6��2�����u��]�^(F��,�v��.�H9�E�6�$�����E���Ԫ+��X0@�H��6-چ""�Щ��nv�%r0S%\���%�LM\EUƶ=F�mQ�hǇ58թ1%�Q�a�⚚�X�`ƶ���fHDH��eb��h���b�4���)2G�-��Uk�*�\�2V���DXB3S2��*j�絥5s-���!n�Wlŭ,��;.nhTp,��-1v;Q��tݲ &Ƶ
��+
��b�W]o��2v�vof����Hh��&3Z-`f��`p�tY�79܈kq�n�#ti�Pvh��0UhSp��9�N�X��l.B��[Zs4�0fL�׀[,z�n�u��+������� 8��,�GF�Ѯf�vJ�6X �˭c��Jk���C�k�� ��W.&.���Ĭĺ �����CAm���g˥���,":��FZE"�4u��eI���k����b�����N.�HGߗxm����%�3�#��oWCL*��)�����ě2��2�j�j��	�@�-����%,J�e�E�6kai*��tF�3LRrsG���c����d�Fӭ�!/ll�m#T &&nS5wk	�7�3P�����R��6]���Gb���e)�B̄6���H-�4�s��Ī1zy(4Ս]-��k5�,HZn�e.H6�i]Xb����5���c �tI�n�-]Y�eTȸ��l��\�][V�.Lخs�L��<_<�X�.� H(䆠���4�h���2�A,�;�6;V���"[uh���w��a��@-f�5�M42㪀V�G&�c��i�j-��*d!P/T�\�)�Ɩ��ui3.���ʎ��i��*��F�f��{4�H��0��#`�J��Jvڳa#Ɔq��f�V� ��[0�Ԍ	k6GB��-lmD��S,�fi4��#��֓5�M�j�`�����3͔�^�1�j�\[�cD`�#sw�
�@�u0���3���V��P��JX�� tIS\��0���b�ۦɩY�.&�. � &0��p��`1f��k(bh�*��e��rPi0rн���F�ZACBX�DU����50Zɻ\s!����� ���%	���nu[��r��u��^.�(�]ųg&����^��b��k��`D��[�$����lWY2u!F�n�UuW2ᘅ%��T�vet�-%��\�ƛS�o'��G΃u�X�sl!nfgW���f����7V����*����g��ٙy]��E���ip�� ���h�G12m�Ħ
Җ���b�K13ke(0ʙ4K+Q)����M����hc,��+he���l�а�9*��]��M��=V��\�W4�5��iEt��PhK\���� �٤�h]�Q�J�WhU����_4�*���ceK�� �8��`�ie��V���rˢԻ]���@�s�R"��5h8��WMt]������V٘����T����[T���D4٦���iP��!�5�[g��Jƭ�k�+�ZB+v-�F,ID��Kl�6\�#t͕&�Y�KrD��mZd�җ�H�T�3�ɩhcK)��H�]�m\�l��LDH�]l1u�Bh.Y�e�ȖU�tA6n\ۭ�Qm�Ƨ9Á�;�T�qF`BضVmp�����[r��b���hYv���RZK�JͶ͆�yrLE5�B4"V	����-�3�f R6g8���i��mv��cp�p���IaEq	l�$#���1�*)��)��]��
j�$r&�^��#6ծ�S6��\m��l\���g�]��%�3�ݙ�7,��SWk��:�r�u�|h�ۋ8��TZ��l�\v��,6�-ZX��8��K@`VV�l4ՙV썚�4�4�Fj�ɑ��B����ysx���5t&�0llu�6s�a�`�#�x�J詐6�%��BY���4p��L1e΄�MHtF�ꆰX�z�[Z%��t���A��)�m
�[���R6�10��2�V�@6n��J�Mz㖀Ձ��l��ZP�]�b�l��+6lnf�pL$m"]�H:�6ˉ�]a0"j%��L؉��P
�P���M�[���Q����,`�)��WQReL�sj�p�"Vֶ���J��]Pl����^�Ky1
��۵�h h^i�M++JF�l�ڎ�R2ʵ�x���Z�gMQ�͓Qn΂�k��ˢ٥QV^B�`�B,��Vhbb`[$��&�,{&6�]���]��<�ݥu5TL��& ���j.îV��c�����4 �\GJ�f5e̷ �R[�-�ѵ���-F�V���e��{L��uX���a����866��&�U���vul�`m�%-aK�k,Z$ҰX7m���+�6�Lɢ�Z�QF�#����i[�Ǌ��
,Is�7�9��ut.��Ͱ�dݯ�\���5�i[���]z�c�c͎h
�bZZ�ܳ�l�P,[��i�*B��[�U]ePk4��Ɗ��geX���T�t������?HȪ���Ü���Ý�� /�������B���G��k�T��E���1�2��t��p\/-Uf�u��vK����=�� hy���#v�����\\;=<w��9�zz��gD����Λ��+u�^�{���gǸ+���0��h��N��JE*����U@6ij2�����wo}�<��Mr+����Ȱ�]�����%��+�� \^Z6z���Ï�o�S/�USM�n��=��x�d�v�d���xY'T��̱�j��]C)58��K��l`j.F�tEZ
��[uHh�Õ���9f��g�����^Rz�3��Y�A�Y+nin⡏Tn]&1d�j�4
�{]ξ���1���&g����D�K���:f4��qg4W���o0�f��݋��w���x�*�,���y��&��X�z��w����菩z1웯��������e�=�{	+�ɑ�g�����B�ګ��^D+������+�[���{o��ժ��Q�f$(��Jv��w ŷz_t�c�/
��|��~Cf�6��tY���6�K�ΔW�ix�o���{�'*ap-�W-�\�ok8���18->~�Z�;�x���8h�$�nnЄ4�Y���_!qGou�띗٬e����'k���ζ{��x�{�];ꟻ���yu��� �1���^QP�h�Y'v�^�H�6�E}���7Wn:*�{�xoT������v��%g�����E��rWh�����!=�n$g����<yv�A�>}�¶#Ȯ8߃���o<���yg�{k���wS�~X��O��;���l��~��d�z�5�o��jA�d
O���k���죧��<3E88���=���V����L�1�ˇτ7�x�|����fP}Vk�����m�{Q1�f�q�9d����`�A�:�IAgz�0�Av<MKD��i�W��w{���}a��V�FsԈ�Nwc��y�,��]
O�/g�_px:�B���IE-����̽�N4mNm�f����>~�*�����8	Z_����:���j֭ec՛�3t��(��Ӏ��s�q+5w�4OOr�Eݳ�$W�O>�}��l�0�Tr>�n"�_N\��dѴ ^�6	sб�\�S���aӗ)_�*�Ƒ)�C]�Z�,���Ś��c*i&��w�j4�Z��^of�IM�ۼ0�m��l�<$�ue��ooQ���m0���)�>g�7~�z�9�zw��K<Z������L<��=1����FAo=ݢ��$IH�G1,d��x�<H ���皌��m�z�O0��g��}�F}��p?{�}���ǂXyV[3&L��C�� �xw���vx��K<��#7�}��~�z��yΜ��q�ec��g"�F��Sf�FRŵ1#�mI�c��Q^�^u��ŏ����)��E>�7����V�X!=���q�+=�z}�W93�U�\��2�8ފgZ+�F{;}�I��{-������o�e��͞ɝ�l� �ˈg���妕[#<���m���ˠ:���0{]����a��lv�ĭ<�5���C��{F{�U�ך�x�d�o���o�4!Ƽ���B��>����4�%�0�*�5����˃"o݇�b �� ���ODͱ�\=D^?;�̐�=�\���{Wˮv
/	�p��\�Y8T{��)�|m��m��xg�`z�x XBPvF<�M�Ic<���_��Ǳ�H������f��#����mh�'�])������S���{������tm�
x��S����s�s�j�ѷ|)�x����o����3�����&��pָ]�'u�F� ��R������x+nw7 P(���ﳼ���4�����_�E"�Q-�v��a���Z�zG�9�`��R�=��Y3����Sn��ׯ��h�Pc����uv�����d���g+4G�k�ɗ����,�����K��4dȌ������m�ulf��1f�c�7Ƕ����!t��v[��UK�*ٺ���b��8혗����#�o\.`n�{�-�o�Bx��G{Ӊ�Aˌ5{G����inN��Šj.�5�X��t����sc^%�D�(]�{cJBb$�N�A�E����z{��ƕ<�/B��6�Hg�HUn	���n�a�Sv"f�����^�\%��sJ2=8��]�Ñ,�#�� :�){�yb����}t\D���ʰ��@��ml߬�j4J`<3Z	f��t��  �m���
�:A��`Ղ{{ �g^C����;F�������*aLk�T��W��a��4<�.�	��OA�Ƿ��ؕ��k��z���"���oIH<l'���u�����?�$)=W�^�����8�c!��Z=f�N�y+� g�wҽ�<k}�p�<W�C2�/9.������12e���ɍgH��n\�{=� '~z�ύ7�rQ+�3���yH}��Ò__���8X����M��}&��8�^��@���q�.;��0���k��z?88��ޛ�@��{4u�ɻ$¼Oj�P��r���]y��Yez&����x��g���?+{#A�I�����;�q���峱���F���m�J��ف���0�aK'���q�9������	�,Ғ�W�r���{��,�G<9gF�F&,�l�ػ�(ynA���7H��AY��z阝�dV�x�BC	XN?7�I���[��և9nz͸ ���ؽ	����irfĈ�p�lI�3��W���4�q��J�OL����w��pu����Qr2�޼&Qӽ��8���0��K'"�a��J��[b�^�9���g�����p����ݮ?Gh^���|UZ����F�ت�T���kZ��v�|][3��cG�R���oxQ�>�sr.�����w&��	75�0�0J�Jtxg{5b�-Vhg^����[����Eoxn̥�x�U����F�]�Ƿ�ı�V�:K(Y�.-Ȩ�:� Yچt��z2\�H������T���Rܱ�t��i�ɜ�!Q�YV|�����N�P�*�s|��g��pD��/��ʳ{�c�k֬Р�$�;��*�F��{ޠ��S�O��/z�o�_P>�o�p`>�*���l9��ށ�+��~��ȅ3�B}4S��
K�wx��9�su:��y���_kW�K�o���d@�ru��Ntm8}����}���n��v��]�:�'l�kO���.�aҘ8I��n��w�/O�����������^x��������2�qu��n�mo%��=��4L~�Ə�t�� v�º�넘��\j��
�Xa�<{�Q7�)�i�g'�I���}�=�6�=�w�D�������1���u���B�0ŸR.,��I˱
!���R�'V�1�����7�X����Ow�{��A����>^xg��؏��#�}Q=��x��R��_T/\w�zx;*��$���'�Cټb�!�VP�Xua��h���T��B���i-�5--�B|�p��w6����<�9z�e����D\�xd�1|=s��ǇEy���_���}���-?��"y����=�I����a�^���ē�N�ϠB�����T5�Q�,�l{-�3D��]%��yx�Ҥ�5$5�tg�����D��`҇y�3���ݼ�ۚ�w���z����{��_^	�|�}^r��'�䞯`ӛ{{�'m'��ͅl�[�{0d�"�l�UP���Kl�a�`]����3qn3�fsA�H/�l�Xj�F$7�q��=�<�^3f��R�O�Ó\u=���g�v�L��/�5�r�$Y(ra�K=ApOp��=�Z��o�+�o|3��r�u�;�؇B�y�%~�Y��Ud�aG�w.-SȥkV~۬����f���.�=����r��{,G|�DU�)��ۋ�a���Z�Ƚ�'�OS�%6й���gN�X��R;Ӫp�>���s�\7T��i�__B��3����m-ӪnL��mV��͗:���ь��y�&����^/w���·��^L��l���-�.�0�Ļ�X8p1�.�ew�Oa�=���?7de|�M������������_{�w�b��9�b�rz��0���r\����F�?i��a��;sV2��^�X7���������}��5؟��)�X����K��N_K�:k��7Ϗ��[�2��oJCc��\8��G��q�)�c�����N�ڧG��b���ϯ� �(@ N�z+���z�&^�%>Ĳ�;����=绞6�;�S��6�^�<�Fؚj�Ё�
���h^~w����8�ꞷ�TVG��,�B���J�Pͷ�v$_�y�.C|}Z&�BĖ	��]n���n�y��"o�
J�����|�v8��Te�}���������Q9�6�sG>��߽�Όo�:V�☜U�e8�!N��q�ڔ�,����6�뾹�o��
���ѽ�aIDw�^�}Gp�Z�����N1zh�ｰw���}��J�|t��7Ga&��,��f�4U/*���JRN���둅@�۷�7&'w/��F����B�q�'��Cρ��r�'�vd$|��Pq���׽�S���S�z^q��y�������{:<��7ݾ�,�/>�ʮ�78�a��Xڴ����K��K���z]{{��n��#�.E��u��G�&��ĝ�{yV��1q+m�|f���p{��S�^CZ�<����P6,hzh8y�o��W���⵩��-3�g�C��C>K|~��{M��לK����1ϲ�he�Ķ<�-">��?h1���*�Q�!���,^�8|rqd�joz�y���y3���u��cݹ��Zr�5=�&�.}g���m�����&�I��ұ�-�+8
t(-V�kP���#'o�ة����Sx�V�3gs}��w���JR�͗��]��.z>n�ﵞ\�ɝ��wpI��3d�Xc�l�q��N�|n��gx��f̣02�7�Epw^����F�/�������=3=��UEn+[d���z3����a@��8s�J����nb-��}�p��4�{e�|�ۢ����/�>���� [�-��ܠ���|�ŵ��C����K��ktL��5�<w�`{�#s�oC����=�v}Ÿ5{V-�}�C�6�%�&G��]�����{��{,/T/���u>��K��}}^P��U�o��'���=�M^/���e�:��b��8�n�1�Y:����f�d�ȊS��%��K`fÑ�Q�;�7��|zw�=��ų� WX�,|wkY�e�2i__.Ƶy-�H��,�kZ<���~��Mٛ�b��~�/?������r�'l\1����;s��8{|���K�k,���\�YX&�j��Y��9X�'w&P@���y.�����E�����V^ލ��xtޝ	�x��{���{^���6^G�n;Q̴̓��άm������|��q�H��o��ok]�n��wܹx��k'w��dtwM�x�7�!�=�ۓ)�����o*��t,Yp�譹P�3���܍1;ײ|rχ��op��@��i~���.�6_m���|��*a�&�*�v��=���[�b$jÊ�%m����ؘ*��2��0({�E	:4L��rk�?lX����s�Ͼ�N���W��=�.vs�˹���?6�s�S�����ށs��}���s�>��ZX�)Mk	�}w5|����;�y�a���6Y3��bc"�e��u���BV;�d[�tG��|���/��/I�D:�;�d)�H;^�aֻ��^��WMx�����/����>��2�Ը����;�o�!��)f�j��jd�I�죭d�雼��kaK�;�kpܖ:# s���]����d�Έ_ �{g5�WՖ���������^���oo�7�Gg���+u`�}���>#�zs���'�M����ok��{Ę�2��|�>��!=dFI�'i�j��rDj���3Z�OՒ��ٙ�@�I&�C�����c�����R��ѻ��?jw;�B�S9�03�.^ˍ���=�[��g�'H+�t�`h5��9<��7}���s=�����Pn����2�}���mX�{����f*z��������Ǻ�gf3����'������g�C���~k�Rƙ#b��P��HV��`#hw��m�j�ӄ�Yo������筍k�$�ww���/����հ�ת�5]��l�4[˞��;�K��ަf��zJ{W2;M��9n�f�}��Į��Qr3��ylF�!�]	�0�3e��~���L9ޫY�+�ˮC7U������f{S���W6�w�Ή#f�f�p��.00N� :��d�����Q�w��������*���v�8�Ş��4 ��^[�{���}�｛ٹ� �Iig�@d�{i��e�ԫn2�V�f)���a߽@��B��<���G�� ߮:�Լ�{tއ�}�-�/e�$�: Hx�]��"��揸wY��z�÷�9�����?Z��,'�����:�����|��_���{����:���<=z34������P�A,��K^ȣ�c��Ŏ`8I�.��v�� �r]�E�f�R9�F��6��t%��N(�eR]fɍ�9�]�,�mT��M۠�^�mR�v"�GX�Vk��1�P��d;�q��隹����X�ɪփ���jm��m3"㬣V�].�ak3��M��ghKM��آ7K�%/m"�k�T��Evn��Wf�����icԸ��R��T��Hi�����6�f듞bWV͌
-��0DũhF�Hi��R��WMe�	Eb�:dX���J��J� �m:�e6�j!�YTVm�$���C�MB���\%nf��V��f�M[����,�Q�R�/i���ѕ&[�ɦZ�n�m��󚑸��CF���B�]3���뵔H�-�6	25�h#]1] ��=�MK5�a���R�ź��Y]��-H::锁��kV�Q�6JE�Bdp�aX�)Z�Zmh�����4m�scT��M�p�3E�M���2���.��!�AU�)\y!���P-Ve ��)l�\@msU.��s1�ݭ1���t��6�f��[iv5�36�[+P�E�mqe#n�UyT4��#��#+���oIZ�Z%663SV�j�#��j�ric�a�����ɘڱ�U�:�c����uݨL��D�򀻆d�-a�)\�lKa�AB9�˓i
��1Ev�It�D������	0�Ev�Lh�,ұ�Y���$�ٺj�fZ7b�G\h�165�h k�m]�w�v��X��`����6eYk�l\�=s��b��vkSb��t���ԫ�ٹ[B-�(�&v�E�BgKZ�@�V�&[��۬�A5��j�sXJ��[F��YH�d���M0�Q�2ۛ���U���X������M�����YEĴ�qE͎�\��]���~�)CA�����\E
���FSW��?��j������T�!�Bv�޾�FF8��ޙ=A:��h�3xf�զO�&%0��x����"��Iϸ�pR4���wx̟K&�޹�;s��դf����ubт$<N�*:p��)�[�q��]W��2�*������<q%�#�K�a˄�dDJ�����%��"����m���ڷ fڴM��u����X�c`����$����v�ˢK;�{B2�N�n����"�4<l�����J�8���{�d8>K3q%�$�؃�n�� ��1x�q�!�J��A��_��6_(����iP�a@�����}ܲi�<ψ����/-�-���t]���|���/�M;�95�	���iFS��,�ib{�c�$�i�D5��)@���H��z2.��M������HP��&��%��d@�uv�s�g^%#�G�KT�Ki�wV��ȋ�|�/}����o�i�DA0�;�	�i+�̼�Ġ2^+�W��d���2ztc��!T(���<,�G�a��Ϧ)��N6������]ъ4#����KEy�;��'{$����� Fb����C<s	��:mP�x}��RM�G!�լ5N,�;���Y�ZS�I� �Y9�,4��2�ጺ8`4[2�J�4�����W�8Ir.�0F(��i��,ke�Z,�H���jCk@8��:�`n����Kp���gR��nYul�����Y�0���+hm��m�1eKJ�]\��.��GjS:�
&�楶(�;v7a�U��fk�ɞu�-�j�.��'�JIa�^��W�v�e� �jj ��-8KJ��,�YV4 
>��)r˸���N���*QUx��ռ��
t��D)*����T�7�U�}V�OtT�9�B���m
���o�hJ|�p�_�!3J�Y��M+�����u��G;���< ���$�a���5�}��sK#z�Tf��'�����A��M �.`�	�.7vD�. �빴y�EM#{�*iw��b(.,.͚lC4o+�-!�J�+����Jqt�����u����T��R3��~��q�H��B���mso��URװ�bCNjH�J9�{��g�X_�ȭ�f@}F3��~(���{��H�Wi�3�����f7P3;6{YP�Z��Ϋ�t�oB�����F8�H'�IO�u�D�"��P�{v�M+���f��\>��ݨ�PP&�h�)����"�|��g��Z���Oef�1	�E����>��t���H�m
����ޱn��Q)�2!0�7���ک��v)�7�B���u
t������tn�����sPR�2�"�v���b��D��,��.-�mXP�=�x��4�3hS���8|.�X�@j;��p�8�H��
�o#z�:[�xҤo'Mw�
��h��"M#	�t���U#{�R��#폤��q�#��$�E<�4`�UG��+�tR��BZKK1�9�Ȓ6ґ1�n0��t����!6ӠH[��Z�{ps�� G'��&������[=��@�H[���LK�{��M+k���i����]��=��-R9�Ʀ��m
u��wX��ڏ%PZ,���u4�̉r�|"��:W�)Ҽ]B�.��OI">��	4ٝK.�� ��h�5`A�Ev��6�f�"X\-K3�	0��-3sk#z�:Y�B�����>������.��I�H�ۄ����:
�6�p�M���)R;���Ӹ͡]��M���*J��(M�!�ኚG;����݊}��u
r��驥�p��(a��lR����F�
t�v�UD�3�bD��9�S��$I�]I�0���J��[�9�_k�ri���ی�U.3��p�D'΁ͻ�arՅ��/���5��H�!B�Z��o�|���^i�"L�H�ۊ�F�D�]�	^V��͎�**�t�G�v�HI8Q��[5R�B�F�A�1��� MKlա&u�l%ۆ�4\$��	�Q��UB�ff5��������Z�0a2�8p�&54�P����ޱSK#z�:[�B������,�*M�%7SK�tUR7�%� S7���j��fLh�H"�M4Ä*k���ޱn�wUUݙ�Ϻ*c3`H�*!�NMD �_mMpf��J"������
c*��g>�辞��K͎�O���&2�#�%����^�	6�v��x���$�?s����{��jN�6���U��\8�%$B�l��n�:gKZ��*�e]��0�e��KF��٘Ph�ٵ�!���ɥ�a&��*%[jn�;ea�lƀ��v�$�6y�e!p:�^EQU�u�б���R,E�MƧ3jm
��� ����%h[[K��X�藲P!�ͦ��#a�Ѵ,�еe���e�0Ie΋�`c\�Z�m�N<�l[�<��,�*B���/�{S��kl�á���(�;�\"�n������U]sC"��m���6����8-����f5n���<>�����54���2�$S`�&�*J��
�q�b�7�D�ܞ�鈴���o�	���8��Α3��z>����6�,�2�+�p�Ba4�&)֏���t�wUM-y�U\�3���,k��b,��p�M��Y�tҥ� ́UJ�6�:Y�B���uA�0O(	!	 �؈�<U��{\�e��] �+�.�V�7�K��2N��=誤w6�M#y:{�վ�<iR�P�l(I���S�q�B�ݖ���.�V2�N鮌�,��_K��\L���R_d���ĵ�P��-f�X��D�L����D�3�d��c����	�����{~;���><�������K�̼O���*��Z�b�����֜�&�6W�b����4�T�� -��2�3hS�o�B�b��fD6*k���w]�.{�UH�m
��q��.ik�aG"�0�a7�LҤU�	r������ou
�Gve�� ��NXL%��A��&�֖+��k��H n�1��Q�zڭ���i\S0*ۋ�G��TҸ͡N��<>���T��R�C��i���LR���+��\_G��l\���>ilv�8�	�ÆȈN�wC�*)^j7���e�J�,d�0�<�b�Eͬ��U�W�GV$��Ӝ�v#˸ôb���YU�N�W]]|�9�D��J�}!�8{����7">�@�	$�@��V���fu
�X�ˀZ.
)7��:��z.�ޡSK1m
U�}��u��.َ�	|�ɶ�P�4��*]�÷�]�=�%��yT��>ԣ�D\�\0�M�X�l�5��.٢��h]I�Y�]M)q�F���!4a�skuu
T�T�H��C��뵚�bc�x!-1%��5SCu��|�y�����1��j�������$S���w!U�f8 )no]P��1��f�&��-���A�n��U�vD��.�>�TM
Q;�o`��{���Akp�Ӂӑ���+�j����h�Y��q[�3 ��x
H>���2���+���������0�	 �8b� �s.������N
�m(��R��T�|#;�\�Y�LJ9yB������~�1���jͻ�I�)�U��R�Sl9vJ���0*HE\��n�v�Ck��?G��}N�W��M+ŵ�|�}�B��o����D4������L�m�1���V���}��yǘ,�I�CM
��o�Y����>�}鑓���x�稅��
/�7;��uoR��$��<�x���O��;�ݞ suI9y�s#:T�:�ޞ{	۱H\�=�C��]�q�i�p&��C����M��#EÌc��{���N��P�eB��S1f'*����;�V�Ci�҈��uMT��$4k6y�[5��*�errgKmvH@m�#3C[vnIEv(�-u�Uĳdf�C%�ٛ
�5��YE�qF�U����L����Uêf�\f痘C�SQRXk��bY�2���f�b�R2�]t1ͫE[*mtխұ�2��1��*��M��-tЬh2^`�6�F��J�v�~���o�OM��-!ԁ���������
u@̩�\e�.�hh�w��0��s�ջ5	RP�L��7��$խ/j��UB�dL�,�
LӄiUA����in��UǺD��ݡ]��t�<�A�Bf	��gLȬ�;�	nꩃ���E��0!2�i��]���)�wH�y�3�}�/3kp
N")2���Nf&t�sh:�սJ��ȗ��[9w��Ap��-�-Ձ�D��3^ʬ��)���\�k]��`k��Ś�*"m�����~������̑��:;�I����8aBpYh���F���wY�Ru�`���yv�<17}*�%^��}d�ڣ��Y7Zr:�*"��s��p�4�Tpw���+�],��+z�1X4E�����$�p"@��Y?@0��k�dI�[� "{7���@j>I�ḩ��3�uW| �{z��-��J����P��	!+�+��Qںbb�fg��{�*c5�\�P�.	��*[�S1��u���35����������k.�f�`�+"KL�Zd%RY�A�qi]4Է��G�������̑'�wW}����Y��a�D�Rm�Q	���o��U�Г۽"M���	��H�(0[nCI����ʪ76f~���t,��P�V��"�;�ʬ��p˷֧|�z�˼
��Nh���v]���f�������>�+CW�w�����J��,����a�^��\!q�yL��+�zl��Wf����8o�?Pwt��sX��t@&�������UW�8ºt�vf�Q�	����AX���7�[���f�o�\=�i�	��$>�v�/c���[,��{�iBa(p"c�a6�FG���]͊p�c���E��w�3�b�I����/.N$-���}oX��uF������.�h��N���x!nte�{pg��{=VE����\���XF��X�C5V�������m9%ɒ_a�+��;�{�1ek�����͗ٹ�=���֬�|*�`�u��;�H_q�T�l�ni�ɁU3P1X�8��w`�$�eXN�U���*;�sy�P�|�UWE��B^����=՘�Z®0��e��k8��%�/[&W��~���x�'�L�gpCqwu�:�@�J���N�ǲV�ox;��m�����nne:�Ugl3�&dS�q�����Q><�`3����{�r���[�k����+����=Jw�����������U�:;�llF��V����/x�Ҹ7�OK�m���+臤8�'P�ݧ��~hv�}�.+��Z2���->����E�7�Ȫ�g�Ol��Gq�4PZ^�^�Ѿ_x#:*�y��#i�х�)mW��@�ڭ�tk~L鸦�K]��n(��話�i�q��j�ɴ�2t����lJ\�9���0��p��f�32��B��[*d1���u%�=0(�Maĭ7if�宱��x1������橷�ψ�[��ů[���	 F�<�gL�c��O�x1��>𵾃45���o����[�a�9 ��Vб��[�-����3p��k�Z��v�g�':65�[X��wY�vӴ�ނ�xS�u�8GB����,U����m�5�Q�M����b�:�NqW<晞�ɝ=�I#�t��"tNa�>o��{]܇q�u�wy�y��RcI�)5cp�jC���?{-\�5�))׺7Xڸ�,f�b�k�yf���r��F�>QV��<s`u�ݛ���w6|tƔ�;�#�-�
4��)$7g�E�U��ɣ�ٚ��!۹@�3�Y��D�QBrb	d����@k����K�_B����Ö�<$��r��Kl����P�P�X����H�{�;��ɥ���[�냗A}��,3��Y�Nމ����.�w�\�н��q�X񚇤��w~[t�W}�`����x���:Ri	��gN�x��3�����q�.�W `k{�q����(����{A�;sz䘈{��w�R��������&@KC���m���h���s]�ʎ�P}���o5�1�{��f\ҹg��;�������}�;G�{�ɸ����6��3��wx�?A�w�`�	��!Ñ��(��Wt����$��.m�������!Y��3���o���&��Q�M�V��h�F���&҄s�(��"�-u3��Cfm�5���Íc\>�!���ͼ� �>���m�5��m��5@��w���Y-Qކ���1	�0����#�~��eBЁ�u��F�Q�3����*��᷐�k��}��:��d֤�ֱ�cZ�6T�a�����<�`}���*;�_v�sm@1���9B����I�C:���&5���� ��޽�f��'� ?w>�H����1�=�qۊ��OgL�n�����B�T.g~�=���� ٵ\݇���+7ۇY��M�����.���_���Z ���5�٬�������������}�IÆ�6D7"��@�=6����wנ*'����PO����^��;���}}jhrj�t�
�RiR�����GM���	�c��ʤa�J�����1�n������1]�;� ��{V�X*!���m���b�dɭ3Ƶ3��kF��q
����՛�A��z9@>��6�)�g������w���̼k3�kֱ��Z���]�7���%�A�� ��/;��I\g����(���v��������7xڒ���C��3����A��LX/Ɖ�c9֍����?w�4r#�j=���f{��Q�T����C�s~�>������ċ�D����������_��:Y�<����c[��`��#xL]8�ھ��G����s2��GV�:��z0%�t���c�m�\%�sk� ]$�6[N��;�ۑ�(:6fib�k���ݠ�c���al��p�)�k����rk��3��]5l%�]eH��:��0�4Iv��1y�&�Z�L�9uX`����	i��(7CmE���64)�1�{c#��ʚ�3��"f��(��Mk�:���n뙳�	|�[�i�Q�i�Mm_��"l�җ���N�'��Ԇ1_vf;���4#& �+��6��"㰚m�@Ɣ��B�,G8 ���A�9�.��q�3����Q�*q�#��"�����A�#�?"=]�c:��I�G��������v�b7z����qW{퍫�5���pQ,��p�Iȣ��o�B~�>�3��;��>��]
���j�����dG��~��6҈i1?Y���]cg�3
����Cq�5��h�Q�*>��}����5������d�a$�'�$Y���"7�09Ǒ�-H{����~���;wEn�X���,����#�|��+��0�6t6m��35�B�Q�R��ZL�l�YXJ��m),BaC	�i�D�0�@�ޱ"��EM}�z��D���Օ����� r���SF!�D8b@���������ޭ�g^a�pw.o3����.#g�����N���w��6z����ު:mV��y3�H�t��}p�XyNe\����mۓl�5CE��.���ɍb��k�9����KCx*#���1��1	��n~����U,���o����Q��\���S)"[$�Z��^� �}wt�-�
�^?u�������[�<�A�!2�iA��\j��{����s`�����{^�4Q����`Q�Q���y��M���"�M������Q�-,�^G5-��.�-������g��=�b~~�~��Ȑ��w�4r"f}�V�D�D��~��DQ���(�p[%7�N~�rD���h�,Q��ZD�3���6�� f���j�w��1�/�IB�"�~����~B v����AJ�`^� ��\������EӅ��2�_\��#��"zٍq8(t����>B�;�-],s�e����.r@�� ����}((E�n�5��|W�~|�����ʾ��!$	?F^���0�h��$��e*�0�=׮�����wW{j�D��ᣑ�R�{��o�*��{3�f�g8Ή4kY6��#�b��m�r5T���d�y1��sO"r�g���9��wo����;#4�׭ı�,���;4-�l�ŋT�9V��Cj�l�y�1<J ��|ٯ|ĝ�����&a���m������Z�GP��w����Ozo��9&s�Mc��G�3��4�X�Z��=��w
���~�j���g�� }da�H�����be�0�O�d[�z�]�g�DgW���Z�C�n=�e��������T9;��<~d���6g���{>��z�~��P�q�]j<�GPż��dI��3�=���_����i����nVA��I�<Z�'��VLނ�Ѻ�VԊ���1�);��-���ϯ<�z~^}�s�%��GX��$�!!�!���{�l���j:#�ܫ�,�J!���g�?Y��K�!��X?{��?C��:�s�eFH�#y����d!��˼-z��ɍ֝Twv�e%K7j�,.*�-�iWT�s���I
fX!��LBq�(�?25w�c������*5
�>��6X�J�I�߿<��w�bo��~�`�8�]����fg뽕-!��כ�o#���~�FډQ�>�}�D�"��GQ�{�����SX��0I�l��5v�so#ș���i�T�Tu}�j�n<�gط�"��~��X���,3�	81�?r:��Du�����J��z��D�Lw���9@������&#���k��d�d���Lc;j%D�{��M�İ`�}~��GQ�:��WFڎ�j}�Qʏ!Q�<��R��8��:��sC�6b&k����cSn��~���s��	�jL���X�w�º�SgoD��^�vQ7�Sh��ͩ*"��_L>
���ΩV�4n��J�C#e�b�@jMWb7]5� �éf�ٷ-4J�H�̑U��a+h�Rhk�6������Û(8H1U�*����ˑ`�e+Q-���*CGJ����;T͊+���aV�j]���R^e,z�-vr�lԖ��4�X��Ύ�(��V�6�\�I��j��K33�a��5��Zw�)Šd��j���XZ��8�6z޳���l]+�Q�j��-X1vsh/4ki��\M�hTsO�wo<.����8Jm��n7~�(����c�s�mG��j>�G���?C��c�tV�G�^��5�cZ�5��M�£��k�U�B�r��3Gs�mCq�j?w�NF�"-B��F��ʅeCh���ȣ���~��Q�Tu{��mC���}Ǿ�*9�#�{��j�CQ��c�u�X��s��ZѲ��T�"nׯ�o��j��Ѣ�P���o�o!Ȗ>�����g�G�F�@3L��N��,gZ6��!��ڽ�a��X7���oa���>�Ѳ��T�>�}Fچ�Z������~�[��1�Ģ�塭k�M!(�6���g5z��I9|�Lb�.qn�gϞ�C�\�P�j����Q�Tu{��e��Q��}�9Ñ�>�$�JBb""b~���g���"�'�"E����W��r�q�2Tc�TL�rq����wӎ��J픣"�������K&�W�L���;Ȗa0���+#�����c�Bk0	��[w	��l�%��C�/=���ơ���F��B��c�s�mB� %G�n=ϱS�k$�u�cƳ���Tu_���F����ᣑ̵`���׾6�F���7w�i�=����˯͚iUK�;�<;���7wF��D�>���ډP�}�sI�r�Pϻ���9��f��4�P�ε�k8ƍ��bf�}FډP̰b����n����mCq����h�y0�<��~��Rl��	cK��=l&��*#"h]�6��c-��M_7�����y߇O�f7w��B��c��j�CQ�u�E�D����ר�P�j�ww��f��$�'�"��E����O�}���E����h��*:�;|�����5{��g}�	�w����}��W�n5�j�CQ���G#�r:�{�Ѷ��.���O�W������[3њ+M�h���t��A�^H�n+J���s`��;�hY�	&�a�/'��*�F�^�B(\�ؒ����������Ŧ�Yam��C���}�]h�Q�*:��WFچ�P�}�~Oj]��l�'����t;����smC�3��D�sw���n<����'~�������s�� ]ށ�S֍�F���7�h�Q�*:��{���ߡ��F���Q�Tu}�zm�p�gO�;�'��]FU"�k�M4�J5u*�ūccC�/WQ,���]�1ϩ:9����kSY1���Q�L���Ѷ���5�\4r9�#�w��,	}��n:�ߘ�g�"�̍�G�F)�Pi5؟��CQ��F��D��;�;usmC��j7wF��B��c��j�T��D��]�
���l0��*߼�bœQ�j:Ͻ�*<�,E�;�}������d{ޱwH�{�BJ0�p�0��Q*������J�#�cݽ7̦b�ğ� ���~ŬD#�N{����p_U��Bj�����O�y� �5�?:���u����'Z�Q��9a��N�f�W43(��]냏���DH���[ZZ���v[k:ֶE�f�qM�bb$���^���*�|Mxᕰ�4�!��(���}����~��E���Q���ݾ\�Q*��Û��w|�%�gڶĬ�69%T6���W�(��-��m8��7EX/���k<�ALE��9��7�{�٣q�L���j%C1�o�ɲ�"'!Q�>����4F�{�
��l��hH���"��g��/��n�'!���ק��y����C�D���Ae��R��m�g��%C1�oדi�r9�w^�چ�j�wF��"fv�����s���g:Ʊ�cY6��%��~��Ty��f��13
��mD�xR#��W����v'���%�mi�U��>w�'{���"fZ�~���~��3�ᤢ(�����G�?�����[�^���O~X�e)��D����8�r��Cb���h��X<k*r-}���7�����V�k��jY��R��$go��x�GmM�8)9���P���C�o3F���H��(��쇮g��_d�Z�[xyG�ܠ���oj��I'���xq�׹X��ؠ�=�݉X�U:�����o�լ�%�a�>{rx�4l�������Z�������� ��v]�Icqn'��5�#0�kY�W������~{R&T��LzJ�t^�9^|�J�֐ă/Y�|��x���=7��_�Q�/9M�K�{�ՄI�yT��r3y/L�P�X�;�h`���:Z{ �z���'�W�G�60����r�NJ�����U�K�@}��q�(�qlI����v�3����k^��;�Ӂ�X}b�	�=u�a�F�K�
jtD�W��ë��z��R)��+��z^���g-��]����Ǟ���ỾLm��{}�p�6d��W�>sox�o<���xo���rM��>�'c�P�Yj���b7���dQc�.�;�:84���Q�3�h6d�d��[ڒ�r���FMWC�\�������1�v�K�՜`����(�{g���ʗ�n)�g;Kk5�DK԰F�$�63b�R3�V��Lq�l��3W�U�����񞺷vv*wfRUs��Ղ����׹�Lj mT;Y��s)d5*-dbVG�b�r��u^_RҮ�xf�����fdG}��6j�nln�sZe�̒x,�J=L#c���]lK�8��hKn��X8V���W��Ԯ�E X�m���D�խu[���C�kL��?�[[�*��B��W+K+
k�8���m)Q�� 1�3�X�j���R(	������Vb��.��I���.Ɖ��lX��%�X!	�q qeݰ���qt�QhG4���B�3g)M���͌KMW�ٖ�k�h6V¶�y�����Ħ˚"A�,�щ�nu+�e�L���%�B&��&��iM5�k@Q��3{Ɇ1B�a�)4͂S��p��l�1Ɉ�K���R#��^UZB�kcuk4/`��v�.pLS:h��SM�l[CC��h2aqj��4�p���5��n�(L�2���M��R8z�CJ�P�l�8 �m�@�u �J��U��[r��|���/�A0ڴ6KP\V�ի,�R�V�Vs5E��9J+n5��.�#�30p�B�"┳F����D�G!�,.�B�w ��i)�ZX1�8��H��Q5rM�3�6,�ؓlhL���G�M �5�tX[��W\�]��MM��(�XrWy�e�(X�(�hl���V�G$%q��Kl�X�,�86�+Sh�Y��In���S�[j�T�%��MM7&�;m�K�q.ĚP*@R��DG��<˚���m+�p�&����B����0ـty���hm��Q�d�4�6��e�G�m�Θ��c��R�c,���5���f�o ��+[�͖��c5�I�2
�:�j����C��)mu����1�vm0\beBb\�vq	f]EHX[z�A�*�F��!�W`�s
;�a�]5a���UTr�ƣ����iE�eu�+v���������\4#G�2ˍ�5	�9�������a#��#PHB�/cS`�����6n�)�9�k��4�e���bÉR����ع�W�4e�� ���f�.���{�3���oǧ���<���ZS�7"���K�fP���$aֳY��,�P�{q�#\V���q��\�4�� nG�ʈ�1M��0ڄT�{��1$#��%\0u��pb�z=�)	c��V�n#�<uw�t7
�9���- l���	�ڍ�/��L�~�2b�GK3F�
%Os�v�8���Jw��OBX�z�n����RwKS�������������\�lL���3遅L;�����o?d�	��vف��m ���3���w�}2{�O��@7��� pˬa�+c$X�@q�~��0�!=р��9��Nl[�Y<$��T��a�!¤�o03������}f�3\#�M��n���޸�# �Kwp��o���${���b����Sr]-�7BĴC�v�k5,8���ѯ`�5�x�SŊ��ƾ���D�wv�n0�Lowfq8��w�=>T*��݌xl㾺.���*�M��lk��u"�f��|Nx.�d�-���Hل<^پ��q�Z.M����VY��!��x>�rx��vz�3u�9��ؗ��:���SlY����k�=��8�O^���H�'�8S�$��ސ\��(�aF TՁ�)cL�%LxO��H��Wqf,k�e=������(t>n�
'g����_( ����pf ]��U���R�kwn� ��պ+v�8�-��I�qS��sf�[���*9�.-�Q�e��ݢQ*3R�t�Hkc�0�{r�������ELcG@.aa�ok.�,�rK��,�n�Tpr^c���VƅIZ�#�q���Ks��(��.�S�V���
k0��Z�Z�q/�.	��3L��mdMb��=�m�:����EM�a��Q�xx�냾��'@t �qm���n����$�:L˶�V���M����-6���LŠ�e��gF����FU�1�0����|�0����Y��v��wݺ6�J�c���ɴ�9»�{g�!���.G�3���h�4cֵ�cYζ�J�c�{��VP��z���"}����GQ3�ۣmBՋ�5��������a]��:yg��>����5��{��G�Ո�v��oԗ���?�G�Gv�D0�SF�P�j�0�}��eGQ3��FډP�q���p�,���w���A�>
�B�-�D�~�>D^wX��C2�"7wF��P3�yC��>�[BE��o��!	�j ����]�V0��;FZ�X�U�bn-mT)6��y��t��j �6'�#�!���c�"��}�d�j��,%F��v �|�|�!C$�	&$Q{����UD*��3�,��
�{c�b���05�d���s�z^�QX{;$n�y0!�sL���uA�Ř�t�ё�(�1�$��rs���6�K%��%Ip��E�Y�M�v۠'mj&ֳ�g�u����o�9Psw�FڃP�s�}�CjA���䟟~_�[vޖ�k-��ȝ�n�9����j%����ѡ�9Fw�E���$iP�a�i� D6$T��1S]����羼��+���Z�GB��]��������N&vQ���iyG2� ~��*�A������w�F �3�\���Y�� .�Q6���ш�Bj���]n�.��:67��t�BdHA�!��IChH�H��#9��
��P}�p���a_{�l�`)�!���Pc�"�ȍށ1�[Q�e��(Y�T7��;�9,
���z�6�
�c���hyG0���B�������j��Z%�I� ��(�G��z��d�����C�g�{��'ǒe=_�u.���R����qV�8���p�­��ʨ��dȥP�D��U���:�w�����ň��LD	D 'Y`���p�r:����ַn�pE�c:܎�9e���ͺ��1��FGp���&���ǽݜ���F{���3��:��A����}|4�Wu�l.�A���G#Ș ��ޟ��'q�jL^��cZ��1�d�jn&a�w.�n�"�����ˎ�������c�}�C�r9��z����T���\�r#Q�l��Ŭc�Z�(9f�*ʡ�]*�*ٳ��>:���m���I�f��o��G#�9����
�P�}�p�j���1C��9ǐs�}�g��s4`�u��bg:6r;������RА` }G]�����a�}w��n5����
��]��|L�1��Z�1��[jC1�_!�����r��AR��������=�]m�5���=8h��s���u�Md���]C�z�a�7�~�9A�+�s�mA�s�����܏���N��k����\�`�Ec������b��l�u�j�q��+�WQ��4�q=��@��t�ci�l�֎',�鵤p6γ�6��Klvې@kV��A͌A��b`,�~����a[��CB	���Cs�$�d}��BEps,B>���o�~�c�_!�����
��Pm_����1��ML��c�2���f�Y��\�Z)rh]A�ٕY��]$�X�x7p4Z[����D�O�߾��w�j���C��1߽��"�T9#��(�$|���AEB�M1��7����Q��$
B��w=��T7�w|4r<��W��څ�"t�����<������R�fy;�z�a�v����ȵ���g#��(�w{��}d#���1�W��xщ�k��5`�Po7tl��a�o�6��c�{����,*���v�	?Qsހ�DÆ�L#�~�>Dn��Pj��G�����*9�����dI�������?I";�Ö�Z *���b��RQ���3[���Th�q3}dcf���=.�z۴K,ھG!���ݐ'�b�7�qr\�� S��!����E��A���.մ��`��i���Ƞ���YZ�lʘ��\�Al�e�Ҷ��b�+�.-������w[�Y��Ba�q��-�����(����4VcVe�?����̶.�HG�CKa��d�q�V��`ݵ�9Q�٣����fԗ]�)�6�+����C�.�l�p�h�(�Ywf�b�Kn�J�?��� �mkII�6��Dm�Jm�-sl��I�ٵ���vt�3pK��^�o&�Q�"m^���٥�+LW<K7nۙZ[�cT�c@sF���~gww+���P�n&3��>��u>�(����`T7D�}��'V��:��뢹Y���D��F7��E���@�bA9��.����a�o�6��c�{��ш�T*:�{�nbɬ�[!�	% Y~�>��P�G�#�F���j%�  ��;�^����g�{"O�G٪8*
��O�`�Ċ?I� P�>���~�P�n��s{��r�!jE@>�}Fʎ���r���R��m�g�=���ߖy;��s-�������n?A�]����"/:���G�B?{����D'6\$�,�F^�(�Wh5@èZ̈́u�;5Z����I�9t<ˡTm�����ؗ���OD��Pkw��Gps��F�V*	����k�@���G�Fo�B�Aa�pɄ�"O�G��$Q��[�9�˒{}�z�mt�=R������"0CI��'	����̉���XDJ��K"�)q7g�u�����壞�_Zk7�шg� @'�v���^[��c�Q;#	"�gډ8�8㥵k�6Ӣ$����^}�}6�w�C��1߻�D�wt����s?w۷�vvt�3��w0��Ѷ��3}���r�"��C���a�7�x�᳑���林0і�m��;�;��%;��I"w߷F�����n�F������@,B��]����#wx��Dα1���3�lwD�w��r�h�E/�tl��a�w駐yǽ�!��3���F}���e��+K����C֕�4P���3��1Ѳ��t��y�P�f�Q�g;��C��}�᳑���{�m�5�w~��V �Tu�۽�Cq�>�򨆐."b i�~�>D^	٧�� �G��C��1���*#P~�}�g#bT�C�﬚�qrڲ�Y�{'{&:����<��=�k;�"H\<+$��j7����=�b��9���"8���F�+��zw�n����J3^�R=�77�:A���ɞ�����}��`��]���ޅV0��y����!,�$�+�9 ��me-���2��H�b�B��;|6r;��Vϋ����G�y;�-�2
i$ď��C=����r5������a��6���u�ܸlwG0���ЌAP�!2�&�,������.��X�C�禚�P�}�p���a��~�T9�i"��Lp����Ʊ!s��Yhf�-حT�-�V^�K�j< �D��{:��
L8i�ÈlH��#�G�ޱ \�c���Cc������P��A���H����#�|^*"!�!�l�S�*���4,D�Tuw���C��wپ9A�;��Fڅ�>����|PL��B@�ș��[�H���{�9��@���{uso�j������?"3:$��G�?�fZs2�G���N�WFʎ���]jC1�~�}���#�Px��D��1SYW���Wbi�^�Ɏ�u���y������̓;�[���~�Tk����{���}��Vw����q���9;��$�D��mŗ[�&Vt�XY�6���_�w�������^����ߟ���F���&�Y��w��}�zm����wF��Q�1���F������GPs]�<\Ɍ�%�F��u��U��t����F;�H��I�n�b��ӣcB�[�he�w�;����Ϥ���aYｰ�n!��-`S聑��?DA�r��&DCR>�r�w�K TC��ѳ�C���9G��ll
r�ތf�C��0��DI�o�B~��FgOъ������>�^Ð�j~�ͷ�vee[�g���'��wtI���o�j�;��6�#�V{�l*�B�����6Tw0�z�mь���u�g�s�mA�f>��hyG2Ԉ9��{����7Üu0��6��cw��x�˖xQ�����32�s��z��ї��Ȑ&t!
�^Nb����
��V0rgd�t^	&�(D3g�B��P�sQQ�9�&��&����)jT�/\�0���ՋF?�f�yJ�X��tRL�a
�&-�]t�KI���.�]�#+�Pu�H�jŚ�hBS���t�f��[�[6��3%
�6�AFVˬ���M�a���f.p�L���T����h�Dԉ+�]��sJj�m1sB�,M�h��y��4Ճ��c�f�s��~[�@��S8���!��ڈ�VRTR��":�蠦�y��\�[蹵�A	��e��-�a16�!5nkL�j�Dߙ�<�G���k<£�{>�=��n5���l�w0��z���%aC�8��w|4<�#�z�]��N(q��"���5u	}���n����m�5���Ñ�+=�����o�5&�k8�5��1�����a��Ѷ��3{�4<��
����װ��A�|6r:��y�����e-Y�{'{�'^��;w~�lwD���r�{�{��@,�Dn��'�(�?ot�2@�|SI-lwA���a�rj���Ѳ�����hr�+���p�sC7�cٗVR����6��d��Kq4G�6�2�*b������������������y'͞G��.�s\��{�p�5���4X0�,��=ޫ4~�>��@P�a�$�.(�����b~�gz1z`���\�TA��p��o�^�}��uY7��{�N��ݶ'�^�j�u�;M�1�P��9�Š�녧����������ŀI $�ٺ:�n�\VV�l�r��8��;�2虰.�;��mYrEnۜ���	BD��@������s�}�Cu�c�᳑�"�r��p�3e-ʵ��y�z�>='C���I蜇��#�z��QC���9G�]�&L�s�cX�&u�m7�Ȉ}�]�n!w�᳐LB���m�B��>�u*�\Gp�����n��(�d};�᳑��V"��_�ϡ�3�׃C��aYｰ�n5�/s��,�β��S���q��Qt�2V,u�	-Ů�L\�l^�b�*{��<���F�7g�2�'��߿?��p1�YQ�1����
ESШ���P�G�#|��"" �ت���z4�*�z�a�n!~����b���q�`�P�}�{9ĽcY3���13��H�����ȣ��ޠ����k��Ԛ:���"m����ZW�I�꫎�%N���ݥ�Z2� �q����dr���v2�3cl�FߢFC���7M���1��s�#K������n6SVr��i���Qi��ˣ�A{r:Z_"gr2wmmkh75Z�u�Rpm�m�E���F�ꓛ&7z��,r��H��g{�9����6�}�D�-�[o��3w}�}����<�p`�v�빚VD��5S��v�N�����9��2�_�k�H�����:�aj��wۍv�3�k�úp�JQ���q�V��� =�y򺞪�� �{����p��{�d�NJ!���~��۬��Ie�j+GZ�ž4p]9��q/��&�L�q�"j�nh���3�tO�_l%] �43��;�ɦ[O��pҩ�o�]���Q���3c�69f��pӎ�T��W2�����:�C'�^'}�b弽��[(��x���QZ�'HX�d7"�q�WT+�;K9Ӭtbƪ�픧LX�!������K������>��8�����v��q����ѧ��'k�l>���, Q��%�� �..�^�z���ً&N������z��6j��ro\���w<v�l*u�`��Z��w��$��^���W�|`~���a�zl��=o^��O��t�3���Ix��W�=�E�{�Kpz]�HpvA铪�N.�n�������rnt�j2�#SF��L�A�2�0�p˓�/o\V�99�����D`G�X�P�,�A�q,��N�Mr~��D0��	���A��7�t�-ԡ^��ݵ\�&���d�{|���Y���-�ՙy��g�v�jAB�H� 1���a��O��"]1��d�cKR�1C��'L�n5�-H"Pi&2%an&��"i�jݏ=���5�~�8ol��d|���%�nJ3�g���p̳T|^�s��0�dt�����/�Z�WW� u���Ȍb洇7tb�>�,���a�?��,���7�LA���O�?U��	�S�雨&�����M(��Ռd G��$�B�Ð?l^�W���x)	�^�
�3'j$�����I,�!ذ�ޞ��7 �XZsfuI��&��,܇G���1h M�pbѦ�D���m���6�D~�e�'�Z(P��F䦁�2�o��x�ݡ��y��kR(S�x0�_vn߃`�>�����;��ya��:N1�z�Cq|���*ūI�}|���c���t�[���9�^Rw&�d����sC W�˹�]��v9��0U���&��k��u|tL;�B��M�x�� y�����X ���s}�f��4��� M�E^�[CtY���\�����|����-!;��K�о��
v�� 1f�RkY���ci�ꏹ���ssH�x`Rg�Gh�!��Qq#�Q�a\��ѷu�V�vi�Eq&��pRgftڂ"��rQ@$$� �22	 X�!�o�}�G�{�����"�B�Æ�d�rƿ0 _�tl��a�n��Pj�{���X�MC5��a�9��v�/D$\�i�LH���#{z��d}ḏ��N\�U}=w��7�{�l��?x��-�H��I�&fH^�"�ƫ1��!Qeݺ���[6����5�l2wx2>� �I�r�;�Uz�e�*)�w�O�Y~�>�(�Ab)�2>�(�;�o��"<�_�tl�C����+=���:w���?~3��L���;>I�~�w�T��ޱw����w��T���z�mt�(4p�6`CI�U��������e�]�3)Enl�Y��]�<ȹ^�oa�U�CY��yy���v��wD��ӵl��̋��ˍ���F����ܥo����7ܛZ�?���	4Q�v�;	��۬-����͑E�ڲ����β��&��Q)�\Q�2b�H�h�|��o����>5&2h0��D6.���*i{���}�NN/w�
���U ���q(��)�SbmD��fmM�H8�r.X�;gK[�X���&�͌a���J��z������G� �٢Ѐ �}���>�b�Lc8�1��Xə�kc��~�}��Ŋ'{w�hT1{�j$���Ð�1V����(!��ؚ1��0j�M}'���R�}�]�*�_��l�C���3鉌MjLkZ�&3�hr��#���G��I��!ȅ��᳐F9���I"ۜby�PL�Se@0ّ��G�q��!��@o�tl��!������܇�D��wiCJ�uH��uP��qU�S��P�,�	����Y��,�Z�}��m�o}qeԨ����X�RdWq�gQ�'�I�6Be3Bh�s�3y��g�i�6el�vX�s+D:�9�^-���E�*���j䣸�&uYv���f��1L\c�j��͚�af��q+�V5��](�a�-�t���D�j�R�&Ԯo_��V��,&Sc7K��1�鑢	6Ŕ̲��7V�F�H5�A�kf�GYKB̈́6cq�Y��8����;e���IHwEӜ]EQ9Rwq��$Q��h*#�(�����qVu���ӝ��e R5��ɱ4�뫋�r��"�L��x�.����.8mLm������wwr������M�q�l9D>�~6r!�w��Ғ�}��/�}�]�u�g�w�g3XεjgY��E>��ٲр����@�I����*����-H���4cשk:��֍�#_{�6"V;�lu'��Y���ݻ�9G��rg���:5�c����T{���C����D1�ݚCp�9�k����
?����7Ʉ�
"O�wwP��K �ݻ�hT1��wğ^l�DQ��?z����	Æ(L%�1;`�1�]eeb�nɍ���D�.���H�F_1Z*�5��{%;�|���zO	N���f�p�J�o�mH���ww��G{��RA���� '��@o¶v����;���2Os��{��'s0�̪;�&2]lD,��V�ڵ{{�I���"T�e�{��}5Τ��-9��g�g^�t���� B� �&b:q�twvw6ˢ�.��+�Ք��3�뎋l$G'G%%�WwY����®��g"�~��%��3=ޔ��4TCFf����HC?��BN@�b ~���9�7�������t���um+�:z=^�$�I$�~~��ʊ{�Ѡ$�����Y� ��_��?}��Z8J �Ċ?^{~�C�Ĵ	PU�y�D�ﻰ�9���6r!�X�븼��ьfk�.	p�JG�0��/Yn�f����Y�����ܝӻ��yD6�v
�g��;����2M��g���!߻��g��`I����@� ���Ȅ4�_Bj��"���oHrZQR�v�b۾C��k����j�^fLc8��3��J�(�~��P�G� �Ξ2 uuy�W@��q'L۹+�+�y2�c�+���@�+����Ժ7�{��V�=�E+:�d�9ҊyM���������$������& 2!'%�u'pw��pYVQ�I�qq�\fggRtT��GqGtu�ue�u]�bC"�!���dwĞ��a�r$����v>����՞OGw�$;�v'�ۺ6�!���6;�"W���9�j���zE�>�C�"<bi$�l��r�����w��aP�C����Ȇ!ｿM��b6!���5�3ZLSL�m��fVh��Έ�Κ�&Q7n6K�"�'tˈ�d8!2QM� �H�H���^��j!��~�9�+�o�e�J�cw�1�G�FwLx�1��j!�Ȩ���p��h�pu��͵���|v;�#�W���
n?A���\��%��q	�dQ��#7��?Y\3{���X1��c���>�#P{����?2>Df�#W7�6	�����!�G=��c�r9����¡�����D �\E'o+%wMN�\̼�\���������v2D�a썷��YڍR��u���Y��-�����t������������>>�??/yt�DRq�_��㨣�������8�.#�����:���9 J�)C�J8���9�#��$B�$3����1�Vg&}���s�L`����;�}�B��1��Ѳ����shr�+���9��z�~�l�[�����k���!TfB36��%�\����ܓk�{$�f0i���6h��|����a_{��jC1�����Tu{���C��9�o8�/3:ֵ�c1�����.a��M�-B }G��c�r9����¡��w�������"NI�ϟ~Ń�ۛZ9O;�N�F����9����T9T��C��Ѳ��9���smA�f>׷�8��Ѥ� �dH�H��>�͟z�ő���'g#�9�k�g�mB�C���T9��1�6KA��P�I�h�d}��BG#�9�	=۫�~�fv�p�s
�� Y�@������?xO�B߰��yN۷��,usU�9�������X���e�J=A��?E@�
e�ZEM]��g2��a���Ďq��	�|~pJd��6���X�t�����b�[6f�B�e�	 ���ݝ�fh눗#`#Wj�-jg��[���#7:���"&���#�z\�R0�3L�m<�q�F��+2̦��yx��lKy�aIHmL2�Šh��9�u�.�k����U+��ME˫Gg�F3A!V���iD�M��1[��%�̔���Eҥ۬��ld'� ���aŕgrD]�fwq�ٝY�q'q��ggE���\q$w�m�m�@$��m��\�7b�,a,p�WV1��i�RkH�ƦR�2WTЖ;��/�0�p��1�kSg#���v�smA�f>����9���o��Q�N��o������� � �8 �f~�>��;���AR�Q�>��F�߯��9��+�s�mBŊ'��}���39��O�MBNG�E��ސ,�?Yޡ"��`�P�n�m�C1��!��O>_�Ի�-պkWΞȝ��gwO����Q����.m�T3{�����G?{װ�<�A�Ix��;ֱ���&��M��;���jFш�n��y�v�aQ*���m1���b�X�ik�4���[*����3ř�q�1v��3h�g"$��;���>4�4��w͝�z}���;��Uw��TJ�>�l��r"7��3��������Cd�M��'􏤊?"/_t�f�O����Q%;7��č��+M�0��OTCBz6�gn�ڙ���ҥ���Ƈ:\йtOe����K�,����9�V��nHq�zv�:qA~;N���ä�q8 &�i���n
#�f���,�Ȧ�HF�ce�25�nl�s0���͵�������B��}~�"�N
dD70܁dQ����z��?Qþ�=6�KV*�CQ��:C��3�� Y�d}�I��l�4̊�`X0�;ۿ��A�f7w�!���w�
�#P�`+����Q�öL��0�l-�?YY��_H�H��X�>���CQ����g#�9��{�m�5��3�o�Ěь��@�A��T���6ie�c�l�i�� v�{;�O5��fBR>�,����z@�(�d|~�l�y0���� T�����]�w��v'��>���S1��s�������l�b �����m�5�����9���aP� 
T>��o9�=Bm��I��?G��?����~�ͯ�}'ֽ�:�
�VS��W�v���tqNơ��
��5G.�q�R�-=YVYev�D��B�(≇d��� �ۼ�T�z�<�<�8�>�� ����N�YE\�Gv֜�";3�肎$N�9Bi�8��9�;3�������l*�A��f��0s�?v�6-ݙ�{'{�;����wZ�#���{
�#P~�}�g#���WP���5��s���ѬMbkS9�rc9ӱ�9³��¡��F(!���`�}�Q���3����9;>Γ��}���qU���]��9kA��خ�WE�h���Y�-�a&/�:I��Z�6!'ZN@�(��}��BE�";6���y���vZP^B��}�]�*읾o�naX��fX�<����OϽ�6Ե`(}F��C�r9�>�^¡����p��ڰD7P��ٳS8�LdɍbcѶ��3_���p�s
�}�Cp�H}��M�`�}�P�����~��P�F�m��$�}$Q�X�j9��{����7�g#�9������L��u^�����ݢTE�s�$�L�\J�.�s_si�t�'M�@���w���}�M����6��B��`Ϧ�f�Fa��9%6ܶ�;���δ�>/<�Q I�ݥ���!'$BN�p�8rHZ&$-GwN�p�s���q�Lg��!'#�D�d}�,�P�>��}�݃o�~�cw|���a��}��r5���|�Z�,�ѹ�n�\:8����1f��m�sE)^���ؒ��'xژG�q�i����s�i�C1�~������߶� ���}����G0s{x�1��γ�k85&3�mA�������
����װ�r5������a��O!h1;��{���Ϯ]�L�h;����l�Ϯ�Ơ�����G2� .����o�#�!��SQ~D_l�!�l���bcZ�T9� wں6Tu0����A�3w�������������xw�w��}��S̒�S4�O'��;�{�m�5�D�wZ�G0����P�j'�ϸl�u0��~�o=:M�>˱j*.nX�}gG������UAʝ�D)�5�,�8�7Bk��F�Z�X���o8 ^���7��#o�dV?tPq�H���X��q��t�m�%��8��ǻ����!��˘|(�o�*6�mP3�F�Et�&7�퀞	��yV�'yK�܀�j�KH=}s��YQQ�^��g=�t���a��z�w�9�d�`����e �u�j)�;�{^��6���=pp���]��{�޾-؊[Gt;r�;0/v),kP���>���{#���z�;���Q"��Q�Al�P�7�n+2�uh����E�ӓF �V��Vl.?q��2qDց���_�/ok�};�v�ztR}�\{��&s�b�^������n�O�L2��8�{7��3�f�����b�h���3v�9ձ��t�;�=^]���&�BJ�rI�.��9{t��L����qF|��%H�x�K��ܚ�}cGt=����o��w������l�;3U{c���:�3+zu�.�LL��YsY8�C՝r�JqQ��Ջ*�������P����#���2��H��
%�w�a�S"3/��l�^��#����H��u�Okε�چ�5��b֗Y���]�/��	�͈QnJ2.�2�7R��=��e���y�WS����F`״���8�LL��y��z�=��-�z\1;��_��}����y�~��\bn w�Bsq�׺,gu@�nUß�����"�'(�,��ލřݤGެ�&}���VP#,,лk+1V�;U�k�WՋ�*�%�L��hp`��Hf�X`��`�]��#cr�#a�����A 7��B�@y�%��n�1hLG��&շ�f:&���kT ��b�ش��b%�m ����4X����a�K�=�v�"V�ͳ	a��F3m��;L���CJM�t��$v�z�ԆM
�V�
hg71��3���X�2�U�ѷ1HMm-#V�DFU�v�"v�"b�6����3)��eJ���1��n�(��-sF�U�: f$F�:��j�E�nR�့ mi�������A�7M"� ��hǙm�5��VIie�V���c4�@l�롓�;Ml�G$$q.c�LVW!4�bEl̺��t"Z$N�2�R6����5mb:�k�R4��B��Z���ԺZBdk٥�&�g2�ˤ CV%�q�p[��t4���L�hB�gi���
J�� !���5A�K(�\iYV�jL�J��,G��-�F7Cl�4[�Ř�Mj0Є�
jB�B�UaBZ�IY����]�4HEp8)ث�v�)��-[aE Ľe����,�,8#�	�deS<]��Jq2ڑtf�e�3�Q�q1u�
�,&��C�&�W:���2����f�M(̙;,J�Ҳ�k��Q�K(Y�jT�k[��flvL�\�9u����a63������dk���Mu�L�n -W��G4� �q �,�&�3�/XRX�ݙ�3-�GBU�W,A-���,.���B��޴�yq�`葵�3
��*�$�F�xoi]�[�jd����Ρ.F�m�.�Wq(L��{l4�$֙��e�WlB��)��iJ�6*Q�#-�%���+f`�͋
0�Ԍ�R:�LRI����m��1Qw*	����&{b�k��Sn�	��B�F�v5[��`4w��{�����)Q��Z��V)@4-�*�L�E%5!�L�Ֆ�AS	��,�d�q��M�0"(������-<��wk��.kH��n�����Aw���$�i�T��t�SW�߃�y�����^�g��pgV1}j�d�;Ʀu\���U(QM啉8�ɳ'�v�m�'E4�=�j�����A�%}n	��>�LAqy<��n���ݺ����� 	���%�*>P�m�T!G��9"(V��'��a7d/98��|"��9�_��9���/��x��799'j�c*K���3��*fܴ
���2�(�Ӹ� ���8t=�q��ێ��;\����g<�.�ļ?X���Cc��t�&����nh�6���0�8hը��v�x�sp���C�b׺�:�p��N��.�"8n��z}몰2ɒ1�@BnLiN��S���rD��`�(�O���wy���A���sSLx�4a�:? }�b=r�{_��c;�u���������p�՚`�i�#���.�tk��t�#=�-3�K�x<�x�sf��7g�b�F���py�Fߘಝ`��Yj7hbݸ��NaG	Ȳs
�G�w�`$�C��V�x
�>�n�@�%:)gosyGyj}��n#w<<�k�KN�GL ����n���.k��n�E����PV��[��m���L)aG�n��k�t1��{X)4���ť�2ǵ�1hbn7R���%Dl�v��T2��^�e�Yr��8�#��і ��������ck��K�F-���q����4�B]�ڂ����R�a���4��G3YGBE
�h�e]���7�\� ��U�3B��� pA��qoK8&h��H�m�!p�Y��p�7ϙ�vݡ
�<e��ل��Ye��m̱�� 7s��hB��F�[0�+�ȇl9�q�;���Y�y��3�tL�kF�A�f8����9³�{aP�j{�nl��'�����Ѷ����2a�Pl���G�E�ٽ [�w�p�:
.N�J	��G�}��9A�=�p��<�c���;�*:�{��̽g:�3�LjL�aP�j�|����a^���Q-H�5{��q�1��C��9��O��]��+���rI����|����Py���wG0����j<��;�~�����{;1>?~��4�kPkvM���=���h����o��p�7��H��?F�Ъ�| �=�6�i���2�*0��+��bGS�@���4��)�w/��6���*At�yg��ϗ��w�j<������G03W�zZ�������$�#{{Bd���A��ݑ�j��@ب�}�*�Mt�V��B�{�8n��l���R1Ţ��lY޾�}�5��s'���jT��=d-�ӎ��B��$��ѻ�UPe����N� � � �GƬ�GK**D�9���:�#����^ �%�a���}Üy����9���~ 
8_s�La�$�q�Nc��o�*�8;��w-B�����ߪ��yz��?2>Dk�\P��(,�ֶ��p./��i����z�mD��ﷹ�� �f}w{~�Q=��oY&&��kX����[MD�+�w�j%G�p����LC��mD����͎�bΟ>~�'��;,��F�.�F��;L��n.��0�Ys:�WB��N���kn�p��R���n?A����9��>����Pj�vP�� @��"���f��Z��A��TYΡ5��y0���6Դ`?CQ���!��g�{
��Q;�ss�-jkߡ�O��:Q(����ͷ�׽l�L��~�ﵯ�0u����\�%U�*�e}Z���Nq��~��=�[L~������A��l9M���ɛ�׎�Ʋ�vuEY�QS�Z�mn�ӻ�2�JI1�Xđ��5&������ޢ��l�Dt��d���)�������}�ɵ��QK3��׾ �>�u*�a��X-�Z&P�ثGw�*i{�� >���2�wz�U+�ڧK���h�(B 0H0c���[��lb�c�R:�,hK)�=h����I�k+����N
i��^�W�ݕ�.e�����~ e�=ޡSK7��ay8D�
v��P��U���Kw�ME/gW�����S)�8*!EM#��]խ����>��`˴{�B�����iC&)ݻ����wz��R���n�n�̕��o���~EMV�t'���ݗw�9H�˔���'�OS1L�6T^�Y�6���!C�Gk�I{/��Q�C/�:&h��9�v���	9>&"�|H$w'Y�]��q'A�q%u��\q��U��{�����K=�0�M�,CLR���b�ׇ�/��}�6�WU*[�Rj)p��#��>NЩD*)��u��@�֤ښfP���FPXJ�5LC��r,B.2\8M��]�3(���լ���}C�s��X��^����JiB($���x����|�o\��Y�X���3�>?U>��14bqwukyz�*]��.� #��b��j�In=)�0��L5�����v��fQ�ͻ�����b�.{����dBF!�6.��SK�ٳ�ծީ5���.�_�M���?z��c9�N�M^#w3��<��Ȕc�o*���$tN⃹!�������ᙽYkl�/b4vC��of���q�G�[fB�X�l2LԪ2�5�ж�:h�0)[K���L]��11iXC9�@�8�\֘��D��ieFZ�@�Ŵ⫝̸jiB:��,� �0��ՙ8t5�-�5�bB�1�ܸ]f��k5i��l�Hαy��-7	���jؚ�	�nNk�-ivHT�m�3�v�:�,�p���a�-�c h��M�����V�M�up��z^�YIqGqSެ̋�:�H����m!�<�Q���2��l�r�2;*��T������.��c\�G?{������yl�9�G����ov��{��g}�4���m(�P�N$"!;�k�t�����|����]��z����}���D��ȧB�e�6)R���.��S�}�ᓼ�8�y�Ҫ)fL��0��P0�Up������7H�w���j����Ϸ���k�b"<"a4K�4�LTҼ]�n�>�����\Fo�B�76fc�|0,��"Q�A�n0.�Al�uWVЍ]�J�ӶE�f�Q��_e�Ţa����^�J��u��G;�{���V�W�v�wzR[�M���چm�߮U��S�sfPIB��9��Ӕa�4��:ԓ�O7-�=_P���ȷQ;X�D��{i��Y���w�ʱ���5<׹��V��k�p���'a�#I��j�wz��𰋯���eE�v�Q�E���^<wH�DU�UR=��uk5u
���K��6����Tm��G}�4�Wu�� ,>�zb�o�b��첑�N
�	����Y��ʵ��B�-��w� ����*in���Cp��'v�wuI�����3}��}ޗ0k3jk��h�M|�ʄ��hۣ�5�Yn-���Fhh��c+�j�#������%�i�^�ޱwh�u
�W���>������QK�}��bmC%�I1wh�uW�V�wz�o/P�K{z��|c~<=)���B0LT��^�۵��&��(��:؉�ޅ�On^�m�f�����O�dL�I�9����s�t���9���>f0tvk�xγ�Y����Q��qZ���=�]��~C��3��:�we�;��#͸����F��'����wh�uT�v�14a��Ai:���-�����w�e�9�U5�9��n#��)�0��L5Qy�B�ׇ� ���s��uk5u
T�۾������V.d����f&�Kmİ��j�Uԍ�wR�,�V���<�s.�-���ߞ�1���
�W�����������.�sQ�`��n����M��|>�g;�b�;��Po���W���iDB���Q	�8�z|j�3��{�������43��U��9CED2�^� B�w�m�;�P��z��U�g4̱��b���pMenT���/�*#z29�ɳ[�4"�qܫr�Lk��;NU�����,m*��}�})�r\��Oq����#>#02����8����tGx+3ͮ��Vv�쎳����ޚ5��`�DrP-8ll��=�Ʀ������b�^�J��u��^}��������!tf��p�Ѧ��F���������2�s�^���P�u&���O<�sW��-��&�������ţ�p�Mg��B"&)����������UA�{�5�3�>kw�E y�!��N
i������A�ީ�Z9��ռ�B�+�&�B�l6.�� !���T���U:[�Rj+����~9v������j8I��F�z�{��~�j�o�b����4��r�t���+1��Ev�~̅�G�ɕN+{�S]�nI:b�.��)��D�j�k1��+k�jD3I�Y��������B��`��Y��r��it������X6&^���0�A�e��5lͣW�V�R�!s��b޻[-C�	�����Xۍ4��f0c-�]R��S;D&[5���Jgh���0���3��e*Й�m3��Y�Uɬ4֐�VYYVl��P�G.3WTvB�R@�ħV*��Em0�A,�h��\��m����w�����RJt
I�vw�Ί�B#Z�,�$��l�%��^,���=�Ζc#	n��kE���&�*E��4��&٬\[�1sa
����f
jp�Az��{�ME.��UH�Ο}���[9���Z[���)6K��nwX��cq��4��wV�z�ׇ�Xe��x��PNpRl��>����7��u�G�R���b�מ�����M8fI�3^�|����*׻�&������� C^�x����ҁ`�шm�Ai;����%J��}�݃3�z�M#��wV��~ϯ��B�[�\���vhL�3K�����RŵjYjv��k]�f�+2��S�Z��X��{��M#{�~��2��/P�K�c��	`�
$�b�Ҍ��Q�傹�����u걖��]�4,�yV-�0A�ch\��1��(��+��5[���vo/z�&1k��czh��u����⢓�M��΋$����Y�������츬�Dq�f0��9�31�&&���\�����R�ޱ~}��T"�m�����٩�s��uk5u
^|-���2�����Wˡr*!C�!7�m����c��qK7�b���55��q��̫^��"�
�\Bb�-��v���F��Eͣ��]ծީ5���wDX�
�!�"�F�Xe)]��e����;J:��� Gj����e#��631{��UH�o]լ��=��[��w�]��| �pK�4�l��Gs����/��&��oz�ݮ��^�|.�i�@�`��*˫[��)R�ޱv@��b<d{h�s����W�L�:6n�^�8��u%m)����mYV����,'�	rg��V�FA�o��@O��r����ukl���E��LA�9����=����/��mM�p~�s���y�ЏE�q��7���W,
�-��q��������
���zc-���;jr̞O�[�˯�B0��N�])�~P+�� }_�=���/h�],iʹ��X�X��N��g��N��"^aۂ�ZC\+PscX�()�������+�=�y2�A�� �{sqq���b=$�%:p�כ�$�j��{�4':��7��L��[���O4�B���n �����ߢ+t��c_t�k#�T�;M��\���˾�ǒbh���Q�t�-��܆ #�o3��� ��"�w�1��Y�)��ᾷ��^�'�jK�>z�V4b�0��0nz��r�&���_��#�z����:"��"!���/��!6���n�&��9P��K=��p&��yi1��a�e���nQ`��n��ܻ��9;���Zl�C��n����)�j'0���L}o��;��|�#�xa�����}���<ֈ]�j�ݒp~@_��nxO -	(�'j�Ug����V���
*�ܝ�/l�	y��[�nئ{4��:XGx���<������m���E����kݨ�%aB��t��15w��m|F��U���Q�*'&�+d�p��Ċ�Ǎm��!��`5��<HW�Lr�"�(2!�����UoO�5�Ǝy���5xS+h�{^Ʃ��ƩT�j�=)��S���pL����%駍��ݥ����8A���|Ђ{�:>X���'���wY����F!�Q��腤@��Py�f�����7��_���pf �貘�K��x7#�^��2�j�������u�������rY��X�������"U�BE�����3IY�Jã�Y����~K���ݮ����˱����f��~'q/�Aet�@t��gf�'f�3d8�׀dnƖ���Yċ�ggo`2t9�z��3��t��4x�ŶÜ��|u�Z�Fx���ӾY��Qyp�x��Ӏ��o.�3\6��Dt <p�x2H�{��ͺ�#2"��nt��%��U�uX>��J��i��A�Y�+JH��v.n���!�B�+ ���@����@��~�03YӜw
r��痴����c�Fnn��&��N3L�!�w�D�y��{���<�r���8 �F��a�9 X�3a�q��7벊9�8J��Y�F�A��n��!^T�]vaـ^B�����Y[><�w�5�ѣ ��{��nx痳}YQoŵ���ۍ�PMt�V��s��
S�;f�X�T00����;��Q���;�q�UDtvhu��gv�X ���7oH�s{���������m8)�j+�|y��˵�O�U#��wW��cy�ŪY���!��m��@�u}SK�|]���b�z��R�ޱ������~>�O��1-4��GJhѣ6���&6�*mbRu�Ve>:x�E���eB31~����j�1�����,87ޟ�cw�<�f
j-�	�ծީ5��/w���׽>5T�f�߾ Gא��=-Rl�m
T�����G;��������k��QI^iAp����
b����@}<]J=��.�f�P�Q�a�Nҍػ"�����q.H��YS�͊���-}�:�����Ho�]lU� ������[�y��D��'�����Hvgw�w{uTw�<�Yݡ�^.����8"�}����|����A�Bi�0O�W��������Ѹ���*�c�3+�E��J)c�[�U��%����ۦQ-��d�Kar�Ace���!ˀ���و0Ӝ�[��woX��s�����y�޻v��Ҝ�P�d��QK3hW� _��t��;�뺵���^}6�v=�H3$�1��G}������~�|���rn)n�
�X񡬂�iB��	�t;�Mv�Օkc�B�.��w�����M,�8^eD(p�$�
!;�k��ME/}���v��2��m�Z]۶cմ���_R�}gp�ɒ5���g�K���;8�L�1|� �[�b�P�GR��a�w�nb�x��p�l���:���k�ft�m-G�ʚ�u*@�:�B�WT@�ګ
]�X�..��cWCiH�GJ�X��������ŅuM{�T.�S�Y+����.Ѭ͋���ԅ�5�m-V�`�u�q�!�.ԍ,���.N]R�q
AE�\��+]�僪Ỳ��4�n��`�[%(WpQ��M����Xo�I:�<''���;����,��:����Ӌ$����yu�w1�Kh�ns6�H�M��k�% �Kip�3�1mZ�Pk	��P�0���۾�wiFw?�i^��������QK�Dz"<�e�KB��GO���{}캵�ޡN�v�������F �A����i��4�;޻�]�B���a����]<i���:ID�
��������5w�[��w�]�9�_T׀���{2mwx�"S�M�অM,��v���/?W��G��]լ���x :{�#�e�Q20խ�s���!*ٛ�L�����kiv@J̈H�X�D�Y���[c3�z���q��sk��{��fK����[(�ˆ�iAi3N���nr�w�+��2Y��S�hN�:�p�M��"VJ��pE�	��z�Wl7���n�ʩz�;��޶g�Tk��0H2]�xj`D�OEV����
�n��#��,�Τ��\wQ�gue��\v]x�DY{����~��U���ǖ�k��a�4�-����^�[��.�}�>�W��G�޻�K:))�I�Xp��^��w�fZ;�W�4�7��o�}���UJY�s%!�D$������N���Fw��X�;�)���wk�ᾨ2� ��!6j ���7Z[�]��.���NԲ�73@!	��@I?�m�z�wH����c�������K��<ф�*I�լ������M��{ݣ��}SJ���}��=�nC(a�Cp�M,�z�ݮ��4�z�-��.%�p<-y��Ը0Α�s��������Y\�3'�M����'D�1�Y�=���G�D��*��5"rb-�)Hr]cSt�)93�}�~I���gtu�ʛu�՝G&"H��LN�u��gػ��s>�����A���La�w~�� 5���SK7޿������U��w��3-s��%�b��J��޻�^�]��v��.�i{�x�J<�1�@�&�afҎP�J ��b2Ѧ��-[e�atA1���P�eb�z�U,��v�������9���Z>,@��!D0�H��t���_��f3���SK;޻�]�Ƽ>��Q��Dy(�l�ػ����Ӥo����}�c�b�w��*���0y8. �a�I�S^|�}�̵��Y��.� s仒�����k������f��gGC��+WM���Ƌ��gT�2!�2"g&�b3������Ή���E|H��� 	~�c����E,��wggI��1	c	��"��R�����ܙ��)�Rq;����B�/}����G}����Ιr��'%F�b���
LD9�"ʓ
�f% [cL�4����\֑�Y�E���4aAP�N-�����]<i�7���}�Ǽ��S��<Q�1!�`8l]�9�_W��U���r�'MU+�����x|잯D"T���z�����=��v����M-�c�`�I�[	]������Y�z�ݮ��4�� �=�̫J=���P�,8LS���b�׀�7޿�m�˕�8j�@Q������s�M\s�o�E���u�٩��B�u�k펽�����+F�ʺG�L9k�"�j���[����8�p�U&+��+z'8"��Ґ�0p�4�l�Z�6�%���4�c&L�ƶ+Q�t�)�Yu�,R�mx�A��iF3QlX^Y�u�m)R%Mp�a̙�+)cX[��*X�ֵ"�\[��kԖh�h�Mal3n�EE�f�������e�j���j�-�i)٦�Ў��	f�,Ř%P�mqF��v�-mFW1�1���i�Lhf.�o�����wIQE{a�k�-��gGvZ]�[h�;^�Y�ޛS�}�v@�E�S��$�R=��W5��]E@��U�Yt&�l�3h��YA���FfύT�ꚋ����\�o�B��xĖ !	�ڀ�T�9�:���x���UKw�b��GO��M�{Ŕ y�	6Ti�խ��
t�;�]�|3�����z��f���0ц$6љ�����fZ�z|i�Q��7W��WzźK���0�80�I�L6.�i{�n��+�|j�foX��Q�(���"
���)�	U��A��B�c;%��j�6�p�uvE̷;�[۴{{�uk#z�:]��<�3�z����(�x�
��M|Swuk��W3��.K���ő�s���Ȯ�wv��{)�r��]d�ev��l+ۓD�r���ݓ
�s��w�6l7��5'�UrH\�D������� G�}$��۱�Yee�}��<�8��I�	�"�ʺQ��ƪ��� M_����
-��0�:���*�󺾯 -loz�Goz����9D�l��M�������H�����oP���~�{e�||J��A,��6����Fo]ͯ|>����[��v�:xӥ�����R�S!ÙU7i�(�LS��V��eB�5��팰Ib��X�d02�f�?���7�z�U.��P{{���Mi�����	��P�BhI�͑��]�S���f�r{�_��B�"�Ǫ3����3�!o�"<�(ɣ�^Ů���bmG��o�ֺ<�R�\�3{���o*.ꦶ�������ݬ"6��Td�<&u��;(tz[݃�'�N�>:~3�> ���0��g/���l��V�߾�?~j���B�/6zi�q	i3U��F�qʼ�T�6�Up��\��t1�&h��J�v�z�U/��{f/G�Ɲ#�2�{����7O�0YF̶L"��.�"\0̨��MM��:��^����ݣ��U�!�]�B���������_���k��T�oBa SdDAI�wk���{��l�z�igH������ﾻ{;�Kl��I�SK9w�ݭޡU����_�]�G�Ɲ.�!�G4RM�!]��|�P��"f߻ꚠ&/=겢���B���C��y��C�����.71R��d�{�V�M�Ŗ�:4N�r��B��@�{��v����X8H�������"c�@&���X۝��SZI�N���s���h��*ifuq��������w��Tnʞ��l�Ԧ��6��y�M:ivI��KU#.����Pٮsi0����,B&�do������ާPs7�}����|j��rG�����Ķ�Tޜ� U���)R��
�Gsk��~���IC.0YF����P���5������ޙ��b�Ep[iت� ^ޡS���F�}wW��7�w4;Y���Q�[)��f�7:x�G�����:���J���*���,���SYѲwfÔ;;h��4������
f�zc#eS�ؑKS��{����Т��F�Yq�?���P��㑟iO$�8D��۹���.�J����r.7,	ӿWm�=FW8<�`>Źm�]�_�D��:�,xN�a}�,�o�9w�{lp�e������3�1�mfƌ��d0���3N죚ꛥ���i�T�\��NӘ��,�����e�}�'���=�sx$��i>��r�9����bP�ź��賦�(�����UK�D��u�������;ƃ�+�teLU�&kte� �P8%�ը�����"��'lVn�Wf�����@`9ge��;Xf�\�=��Zw��F���u��O�Wx'�8&_G��][��y��mj�o���4|����^Μ��sΉn�{)��yw�zY����iEF�Ac؇���)���wgq8�9��;���z�^ɫ��k�;M�</��Yw9d��Y"��]k��kVMݍJ6oс�Vh͍�0�5q��-��qi�}i�}O���;�D��w����Y�N9����w���0�C�^G׋��|�
��yaf�����5V�����cu޴s!�|i"{�����>�3��`&UX��M��tx�v��Ÿ��Ǆ����=jw��DE��N��r�5p[�5���U�;G��\��=��
}��Չ�U�M��1�bʈSv�W�^��g7kW�*T�[j2c&�S04;�ag��<yN>��M�e'{h�VnC����#�j
<!�d �
�K����u�]�m�+�M�&ʌ%�˂�me���%a(��b�n+�Q��F��[s��[e6L;:�)V%���\@C1I��m*/Tb؉!
�e��bԱ6*4���k4�Ws����&r�#n�N�e��ICh�r�q/\�`��L�ū��sYF�3eZ˱.�1f.��e��-�PQ2���ñ�6�L�J��m�k��%��WX�Ѱ�#3�-�p��Z41c� �!*S�t���a�5f�b8�Ա�4���2tbE�s���i��[LC$���:c$��d/� �HZ˄�����k@̵���]th�ei�X]��tX�fa5�ibCm������8� �vƌ���+4`�ډ+s2��mÅ�l^Ul��s�3Kk�6�L�%x��Mf��;T���X@�5	f2T�\��n�/3<cC%LST ���c��[�Km��d��f��P�����i�
2��jEH6��.p7@u �]�ݕ�K]�h��Ѳ�y-�[�GpʭjLv��.CYe%z��u����ol��)4d)��@��%0a�!��&x(�0*��o5��-�6l���,����f�1����l��	��6��0��/	l6��sb�A��,��3�n�1��[,K�ؚ��lҙ� �[CJ1�A
�跘���I�6�\Sg$�S���\�C5�Vg�6�[�lK��uS)��6�	{7m��!�BJ!#�P�S;���nB�ť�m�h�m�s�2�����VƷTpD�f:�l�W�VS$8����Ê��uB��cT� �uEe�qGi���Z����,�+Q�ֈƔeѭ1�4�*h����A��е�i�[��Ƞ�CA4i��5v6ɫ`H!�R��h��&U�e��,�r���4n,�3\�mrR�բMfV�%���p݃9XO���%�'�����=��${�G�C�5���z+�)��It늴�n���oEײ=��CQpb!7�}paRT��N�[�Vv�^͉�	ؚ:�ZO�������L>s���Y�~���r��qd��3�X�C����'�������{p۹Qm-W��j�^M ]V����C�dh���}*}�k�8m�7�?����n�x��CS�F|S��4����ݺ� ?u\�=&��B`\�ʬ^�rx�o�_,��5��Qa�/����"�<e�m��/��ۻ�4A����f��<�پ�<nA�y�sN�'�K�{�m>�>�w��(��~�T�������6�&֜�G�]�t����DܱxQ�����u�fa��cK`�&�]�SF���G��
�
G5�����z����tT}��	�ב��]�6O�˄oDf��\1{������]���M�i'��ޒm�o�$�+�3���{]�B���ݒv���Y��(Ô�_�K���J��:Ȼ;�J�PN���c��al��܈�jh�4~����2wtl��"JX�� r��~�'�7���z��~"�9ĺx_����\���y��W���I��ghThd܀tPF�0�0��f��\3P�RiE1pf"�]ibmZ�����c%A�8�E(Ғ���0T�V�AŶ�����(e�Kb�R7 96�ֵ#MZ�۴3d����MNS���W�2�� #-D��S+h�l�\�ǈ�],���^���y�e������5�fcU��li�eʪ!Vl#,�����j�&Cio�y�;e��Ϟy�rp��l�i<�2�H�@�A�u����p�����#�ŵ�ZVm��h�a�B*j�d�q)6�t�;��uh��
�Y�\|٘�=>4�v��<'��!''wV�:g�|�ݽ����*h^�Ux�{�H���J)6*�}�&b�7i�����Gw�J�Xp��)��w�|�������]գ��*k�|��b����(0�)�-&i�7�뺵� ��
t���U#�����}�ؽ��(N	P��/M�sU���7#��c!n���[����i�M���@��&�+��
�Y�B��FΟ| ��w�ꚃ�CɸeC`�	�q��'ӈ�m��l��QR�zv�J��kxP�q�GGe[N��Ѥ��c��5�ѻ����w�U�/�`c�A �A�D�amj&ۉ�v��A?$�⏦�T�;�뺴sz�x�[y�y����Q$�ݮ�O�T��|>�wާ=�!�Vi�mn 4�W�;��z�7ޡU��*���j�z�{�! G�IC�:�����{��������B���޻�^�S��54�L6�j`�f���st�\酀[jݳkr�4�(:�a��
L��b���z�ݮ��4����e���P�Iv�|�{�҈��&v�wP�}�[;��˫G��4�7�{�������o�[t�v���/7�Rw�k�O����,Ě��>�a�{����͈���d>�YN焆	La���&�*�D�S��וn�;�
~�׷ߛx/(�m;0,��k;���CZm���߿W�X�{jkz"::D2�& ���|{�b�7{�*�c{�׾���޻��1�Ȩ�Km"�6*���LǾ�E��͍��UE��O}>���?����lv.�%MΎ#��e��јE��c�˴Ɣ�k�h�-����SB��h�q���:��U��=��\���UUx���	d��4��Vf����1w�9����]<k�}�����3�o�4�]Z��P�K�z�߾��g}�4�o�wV�z"�)҆JM��������h��.Q��uwb�i�O�nN�Ҩv�<9BF+��A��`Lf���n�m\wf�Rl+��1 랳���q[�Yb�EN�{�ol��'�I�!��]����aZkk4kmn�1m���ߟ�)ҽ>&"�����v�wP���>��d�>�P����b�׾�4��$n�([����
Tq�Ů�a���lL��f.��\�sPh��Q�p�nǈ��߮��F�
t���~�ᙌ�B��	I�!��N�mޡ^}V�{�.�|e�;y�|>���!��pS&)����.��S��7�̛G��4�gB�ACd(�	1w~ 㧍9G�z�do�S������ix���X(CjNi1SKc;��׀�G��.mn��]�:�˕菧�$�dR���^<�gA�Fgrz^�Y��i�ٹ":0�\*kGz9F�ú��FY�a��\�ƨm��N��egL�;nꆌ�cf/�bI���L�D��P�@�¬EqF��,qb��eb�ܸ؎FؓT�e�J��4�,7j;C6�m@�#(����ʹa.X�ج���ո�X�G��� �U�:�m�60�;Be�"�6�Ky���VЗ	�:aK��u�e-!��&NXU�i��3Qjfm�ss�6j��b��]�Km�
���;n�V5Jm���+�
_�;��w�^6$$P��e��δ�B[`�W�瞚��q@���7�#�7�GY�m��Rږ���T�-�g�y��0�1��[�w�S�۽b������][��z�my���`��L&AM1SK3z����4w3n��F��x|&���{�ڈ��&!1wh��T������c>�X���ޱwkX:yJR�I�HlR��q��fU�Gz�:]��.��|�}�4�����PCn �II�ͣ��*i{���]�:�M�e�Z��h���D�ˍ*�q	t2,ؚՌ�(�V7G\�B���j�����*!��H�	��=���G;�T������}����B����G��h��i�л���Ə�͏q�7t�d.j�-I�f���b���B�wr��G
޵�:�^]�*��VʦT��;!�4�uL��w���Kn����$�"	 � @�X���m���m�f�L�0`���]Z�oP�K3hW��kO�<���-13��]�ސ����g�u\y�K��#���b?�8p�ګ� N��t�z�U#{�*k����d���R2��5�b���P���>����{�SQq�������J��H[���V1�ikfdD5[��.���WKD��%�a�w��B��Fw]ͮޡ������X���{�SF	��,��f�#ݽw��c�b�-�2�fP�}V�|��JM��Sysk��T�7�]��7/�ON9O��S[c��|�7f�n\Ll=�K-�+/��2��h}B�E��t��&�ym���{c*Kھ2k>l~'����~�~�𰘼HKİ���y[]��˰�5 ��&"#�b&9��s{����� �E6IaBb�{�ޡU(��
�Y޻~|���wIf�#��BE&.�tt�K����eb��P�K6D̯�h��qۃ8Ե*��-%�Ah��]1��LP0`���,��C(4���w{�uk;�f77��ᙜ|�e��z�%���7	L�լ�����+'�6���4���� *���R�����C����X����Ɵ� [=��eZ��P�Ift!xCj"`�b�����X��w{�]գ��SJ�9�{�W��q~�6)ڵ��"�y�]q��w��JWUXs*�MrK+�A��Ooj�n�Gu�Z��qg��90���>��/����,�fѳ����������Ƚ�}���?�Hkޅ����$��:G{z�{��~�j��G/(T������i�ө��sb�H�r3+cU��-�c�b�RV��Us�.fP�Q�����Rs�{��33�������*��뻏B��>D��i�\Cb&/:}����ͱSKc}빴sz������#��1Z-5ػ�>~�[��^��yz�Ln�fb��N
m8LL��-���.���e������G�Ɯ{:"<O�%�p�-'	ݜ��|۾�{�5�=ꩇg#����X�}>��ϝ�}�q���.�/=���d��{���O��4%C��5Ҫfؙ�ʌwX���!��޳Pm�u�&��;�I��P�N!H���XK	��nє)YU�e�`��\0`�r��X3Pl��JI�3E�����l*�2���ƺ롃V*���JD.Ae2���+�6�J��Y����is�rۨ1�D�	d��	.��beX�+t(ĺ73ToG�4[V�)lCQt%	r�Mt��tK��֪3��*�܆t�Í��]�i�([avN�k}L��n�M��\XHt8�ke�Fy�If,F��l̘nT�mmr�-�F���2]X$:��d3@� �L���hMϣ3gƪ27������뵝ޡUǌ�^��ICpXp2�ޡ^�|*��������TҼޱ~�����-��`$�$���IGF��լ��){ﾷ�B�Q��4�<�,�h&Z'w7��7�w4�{�.�lt�^ =�YV�o���[pK&)R͑3+��b�����sh��T��t��C��!�ͱ��4�����n��;(�Hu��(1��I]��F!�()1�����N�׻���j� v��L�ךe�A���Ai��Y�]�	�YfD�q���Q�"�k'���r��&�8�-�gv*}�.�d��A�y�9\��f���[�Ux+�����.����:��L@ �#1��m�[;�Knm<x�~�wUM+��v�:xׇ�m�����m���2��lw�S���*�>���4�7޻�\��RBdi��������k���H���u~�|�w�[��|������I��Q]�9�B�����ٓ���B������^��{����,��`jM3b��R�5�b�qh2+�7�Xdj:iWhc �h�4	%�m�<����doP�Ksh{�ݳ��*i�"��SM/�%�w6�oP�| �y��v��t���W����>PcȔ�-CP��:]�B���zdmfx���P�#������J�+Η�z�k�'u���uGN���EUn�:�X���Z�B�9�[��`�u^�J��.�}��#�Gc,Xh�K���Z-�0���Jq�h��X�
<]\e:��zp�7�٢�q�
|##�4-��ҙ.�sG;��yծ����8_�j*ŻX�+Y��4���},[��]\��<��wO�B"��X�;p
j^�C}�.>� t�������b��%����m{�����ѯ�����=���r��ؓ��>��{']�?v�V��j8�NV�3&��u�+l�ܲ"n�X٥��0#зR�쎪y�뻀C����_v��6�L��q�XR�����Gj0�K]�(9��C[D�E����D�%{����\:Y2�������S�6��)�}W}}f��Չ��W]!3�W;̌Sٶ�.�ZK/j*�v�T<� ���u�V872��76��if����~]����ȸ���{}����>�fڡU���]p
u��}����ݧ�!=��.��Z�F���v�c�D��(�����6T�4\�F�3T��h�٧|Wt�ӱɗ���]�6g������K��d!�7����ӄ�f��1ܔ�oj�u��ۛ��B,�P�I
vU4��p�=���/�'w=�g�R}wy�j��Nq�hَ~>��{���^F�y�i%,��������;� �����5��5�'�+��9O�yf��uZ G�����7���S��퍣]!;h�n�*��؃{f3EY�� ���]8.�X�	���Y����0�<M��#�9�����uǮ�I|F�����{�罨���G3�^�8f�g���K4�N�Ou[��B���'B���q����<.�{<����/��t�C�I���p3��n�ϥN��_on�V�0���3oD��k��;0��>pXXB������A�-\,�����yF:���w����X��7a�O{x���2O����֨Z��K
�	��fA��R��jm��͐��n��yR��i:�[1 ��_�|9��V)�t<
f��0r�&Ե*���DD�u����z���vxL:��4nM��X`[$�ҔЏ�Į��o#�Z_f���������4ȳY©,������HoՏ4�7|;�}͂��_-0~^�7�f��ݥ�Q�;1��67I�9���a>�2���~�聤��b��R\�9"T$vnIw��0�p�O��_�p�>�#�����|��)�^!�5H;tk�::|���{"��,������#%�#ޟG�~+�;�����Ԛ�U���C��@��n��6�'[E��3R����?|��}وt"t����l�n�y��qgh�����G��T��tA��1a��)�w~ ���H���w�K�|>y�b���zS	8ʈD�b���{��ׇ�G��.mgq���]<i����#�v��rcL��mE�d��Wdk��Vjl�
&���n �8u����~z�G�"\���v�{�{��տF��sk��� �d�C@�ة�y�b���1�=^4���Eգ�"|>�i���Ŷ!4[��&�ݣ��
�]�w>c>�X���ޱwh��E80L�d�Х^��=�gѕh�H�*�6����c0��6�$$�ȫ����+�q��l~���$}�����N}�R���)�
9K���t����"Z�<ڽ��+V���f�gϦ�f	����kvY��o�e1 -�B���'�=o�_�Հ��&�7w6�oP���������t����~���}��y�13]360Z��H�EfKA��hd]�c3���z��U�j�U����X��s��M.�޿���w�T�[��!#�������ƽ��m����G�"\������>�I,�a� 4�����z�mޡS���w{]�G�Ɲ.���d�ӄ�&!�W��;�)��ޱwh纅M{�~[�fM�>�J`�A��L�1SJ�z�ݯ����ݣ��X��w�K�����g�_]��\Ÿ�_1CX�gq���ۍT�8����O-�=��*E>�X1����2�NlЎsF	Tc�c�Ե�
�L�#�����]��oy��]4�u�����X	Mf�S�F��.��n�	���`B�$٫��"�Ep��l�-���Qܦ��1���#�l��3u��1j3MJU�shj╄n���5�l�ْ��ZZ�3�¦[cP�hb#3��k�2�9�mr��@2CW4�[XSj]5�.£^"�tq4�S&��u�yLS��� ��1��N�נ�Łm�R�
_=�z�PPdf�u�&df��@��Gh�Plvn����hM�n�J��hp\��~�{��4�3��mޡ� .����U-`��Q�Q"!�I-�N��wX�|>�g�B\���v�{�W���.E��5I%2�����K�W�*�}���Wt��ޱuh��9�����|{���h�U4�7��o�|{�)�����4��a�B��ǧ�:^�{V#ޑ.Un틻]���པ�
�m�-�	�#Gj�\�(T��fq+Gb���	@��I���L7sk��]ݣ�"\���}UO#Ӧ�.�DG��Ʉ�-����]Z�ޡO��=�:	��QY7{�7�6�f��I���>��İխw6�K�T�+�ͺ/zj�c�F�7�����Vk���O�>	 A!�7D٤��d�o�=|���5H�uT��޻�����Մ &T"�4
hS��"fU�Nz �s��2�lw�S��6�$y�Sl��л� ����oz�����yB�Uǎ�80L�d��f�#}��uk�}��bݬ��UR7�U4��xz�2�M%

0�Bl(��-itсs���2�Y-�
�dvSKvsUw�V#�H�*�D̫�N}�6�wz�ե��ze6�((LS�}�+�}��9�u4�{�wh�H���b��	(��q
v�=>4�!��.�r{�=q�=���O�q�;�8�2^4��\��S�C͉�n�r�LE�{�nhQ�Wo�h�Zt�Vbs/�7 �O� �	I`�^<U⬬��-����>o}]�^��z�U-{�$�Pj!��:���>��fZ=��e�
�����q�Kwމ.�m�K��]Z�ޡN�����T���M,�z��x}��Έ�P���E?�0�<�]�h��<�L4�q��YGl(�Yy��R�ebL���]�B��FΚt��Ǿ�{�*V<�r& '�wh����|[�������
�[�B���]��`��L$�������z�լ��+��O6�L��ꩥ~Q���C��Kn��ޱsK��UR���N���fZc���ֻ*e54���e�'k���9*�˦�6���[' ���NY�gSF�Ml�1Z�q|b4����)���g�8�
�a�J���w�?����J3A^$�@Â�lR��"fW��F��ͭ�z��ޡSK�|��}��ԋ.f"ԫԣCilX�4�R��q̻5C�-%���qC	CLd����s�N���uk5u����q�b��ma@ECnb�����c;ޱSK��*�xg�M?gDG,�����ȵ��B�,�>L�����w����5AE��-�	�S^ �}b��\���*k~���ŪX=ԒE!�8A�v3�fc�}�޻�9Ϗ���P��8T�fl�U���={���i�Ԋ���A�:%TT�t�����={��N�|�k{���A��8r}>�Hsߖs��=�.����V]�vGf�B5�I�����:�����X�r��ے٠��4uG�:����4�L:��&����Z��V��he�һ��E��	�\�9	��\��i��f:Y��L#� ,Yt6�)j�f���RN
�I��Mf.M�����n��K��ջs�H����j�ҕ�m-W2���O�]����8�2;����(�ⷯV�^k���j���Ҳc�P���h�M��Z�1qBZ����f�.i��m�Jp��H���b��j��f�������ک��|כMAm4)Bwuh�O�U��X��y�(�l_ �z���7	��@��*[�B����5<����e�;�񩤯�w0�0��!��.�����Ɯ���b��j�
U��{�b�>�X(5�j	i�SKc��sk�}��nu
�Eg�\���n�P$��n��WB��P��F�G\J����:�Mav�PrXu�ZA�.��h�	%,8���R���*�������z�m{�Z�a��d��Ks�V��ܒ�;g\>u�Awu����Y7��.��13NN�sy3Ֆp�꼪�xS�
�c ��1�ۂ��]�ʥ`��W����"�|$����cQ'u�e������<\^0T��7�B��b�
��|����^%���.��w��SKc���� 1��
q��&b�#��
�O| Q��\�l>"Tf쉞�|��h9���B�p�2I)����}�}���ZZh�]^z߲w����o�7<`�ݓ0����V�У\��+�v�=��Y�n(,6����̦.3�V���U#{�*il{��{����5���LCJC�Zv�~���ʻ4����f�
����\�-2�0�"Sb��G�빴s�Kn缏����e�-�E�\/g�8*n����b�zn�yH��.Ӻ��Х�%Z�g�P#�蟽����Ϙ �β���ͫ+:����_^�
�EwD�]y��d����*+7�|�w�[���*�ݡS]���޻t�y�B-&�p�0��J��*�x}�=�H�:�M+��
t�����(�!�R.�ڬ�����[���s0lj%u��݅�B�����(�N431��T��ͪt���~�T�g�A)�d��4���|&�͡.V{hUR7�B�}�y��~m8-��p�O-�|�8�P�*��Uh [���H�H�)R�XCp�l$�1N� ��]�9�B����S���=�8T�<���
]u�^f��gY��S�Vq�&P�.�^��W�d���y0�7*c�0m�շ����'����ǑqC'�dt����e�Q����m�����.K��~�/_����a$a�C�]�fύT{�gHS�e��$LƏ�Θ1��<��J8*W�g8&�����I���5���Jb��R��Uv�C�%���t{ާPow������U���\Gwxǋ�l4[��]��~|�^抪G=�*il{�������0�)�`� �����ޱwkc��?��s�)�9�%ʷgކ!���.�����}�4�=�]ͣ��*k� �z�s-y��
)�	��0٧H�H�+�|#6�:Y�UH�m
�Z4/��`������p�e�Ȕ����r4����otF%;9�V�/2l��u9/�܎���2�~���g&嗗�C�S��{u��i�B��I�;���Q7q������  :����Ǐp��=�r��@�3�td��](�_�5{<��j�!#_-,�d�q��Gv�7fHΗ�!�����x�Uu���$%����@�������/���ʗ�I�x���i(�辫����2F�P�"��!��?�4�Ƚ�+�g.�,��g���L'o��������S��X/i��彼��ǹ����&��솝���{v;j�}9�%-��b����&�G~9~�w�t~�9.��3nN��TLO��{���d��ݛ�=��QEӎ~��
&��O��ry�In7x��ߡҲw̿�����:n�ݶ"'fɋr�V�VY�g^oJ�Ӱ�k����5Q�u,]nL��yUQj�c�ع�|�w�@�0f��o0�q�e�?���*��Ʈ6v7���6X��P���զ��{�x��F���0
�(��5��
�Y����>��we����.X|]��`|b���0{8,XRc%�k�%�[�X�����0L'�-0-�U^�J��!]�o}��J�
���c���P��v�;�U�Q@�:Q̍S�;{�s:�2;:��韧^I\�z{���W�.aG�^�;�ĳ�nD=ړQPva^_�'ȥ $U�b�P�Ŗ��m�-W0W,����"��Բ��f���`A�C
֩tu!J���n��"��n�B�	������p���^D˪gF�cah�e�c.��(�6��.ee[t��B�#�m��jn�S�^�Ѻ\TR��Xs�v���b%�q.�;�<cY�`���0Ip ��&�R;��]�M���2�n��Y��9�eX�J�:Zf�Q�V�Љ��1Fcr�6.�6ʄh��kKP��Bݦ�SF�����.�к�ɂXCrl��wP���ثei*l��q��D�	�\�� h���L5��ha2$Hh��M5nZlb�!���f1�[��6�QV�Ц����X�6����煮l
*YsN.��@Ø�ZY���!R��g��2Yk��j�V�)�j�@%����jcLj[(����\B�ft�eF�94�#��,�t�sb��*h�0�]nU �+YmP3ۘ.��t#�0��rV\L��Ɓ��qf���+�Y�B���-��sh�Mj��ʔibJ%ljK����\�3k���F�pZ6�\Q=��)
 �T�4Ջ�V�/e�enf�l[�y������>X�!Ǟ6�(1,K,������ƒ8�ɓ/gB+�\�a.�������!�j�Z&����%�+Iy��`��5�]n*�\����`��p�1��Z�6�ͫ�W��bh��NS��F�`��ha-)���Š��4\��p��F�ˁmn�m���W�ҝ��z-5FhMA���Z�V�-0�ݴ[t����[y`:�;�l5�I�����[C0,Ɋ�����R�0���Z�B�����V4��Ba(к�顁hcX�j�l�3vn^:󥱡�f�f![��è��R�����	%��E�tf�a%�7:r�ЩZM-�/�R�ɰ�G��\�vՍ�!�eG6��'�@�_�lI��%�2���K;S�4�"���ަh(2n����my��Մ�_Hp.�M`��eƬZ2�Ɩ��pY�`�W�e�v�&�V9뀣S`�,9�Ӵ@�>��8�͹���dx�A��wp��h�XW���ߩIo�L��'7�X�M?o�s���{�ż����$�;�-��Eⱉּ�?b��:��'Om�r|�ՉQps�8215_�X��QuO{&V��P�p.���ޛ��kE�0{�~3���WcN�!CN��H�IB�a�!ƌ�	GpNr����O����8ќ6�)�hѯF�Tj.-;Ay퀗x2)��}��ymݡ���]�̉P� ��880}��_� wE>�{��R�ƃg~���
b���kl�5b)��5�
�C;SGs�f�W6a��a��5`*ǥf�;���*��{�@��XذN�^9��f�|�s�m���X�]�:�������[��'�
|����{ �n���[��ӓq@���OFM��ݤÓL�j��enM���["������r�ڛ�ɜ:gy���,?w�lG�tb��-�^��i��p���.����p-0� ��|�~�9�����]���Ƙis6]˃L4a�v�t�6�+IlΡA�6��74��EM��c7>x��&�F`	�*�B�K�0��k�¸�X�ܺ�f�T�v�[t�&�.��ր���v	tB%#X��1�8#����cGW`��M�bܦ�B�4���9��g�ƀ56ҭ4����r�}��$�@��%�$+��l�[h賳�md���'���-�!�na�3F��$��A�l�AҥT�7R�`<�鵍1k[$��T�;ޡSJ�k�ݭ��?��smFy	r�'4�D�B%�	
t��B�����4�=�]ͣ��+� *�O T4�L4"7v�=>4�����S9�)��m
�V�p@�RZ�À�M���>|��fM���
�W�\n���/W��]�cșD�pAl�bݣ�"\����v�{�T���u���I�Q�����),�A<��ś$���ս�XLW+lc�P�`��I�W��A�6�p�0�8����ݭ��4�Ρ�}�ճ�"\����\��M�G=�+kvϻ��r�B�q�nMP5Y��E�^ZN7b2=a���R�j"�׵�d؛�}�H�QKw.�1�֜�c_Y|O�T_.�˛wg����싺mvE�Ys�7��eM�}~|���{�*�^oX���{5��4�-�i�;��SJ�6�>�ow�.��SK3���M�j$a;��}�{�X���ޱwk`t�^�|�w�.i,��M�-	�t�=B�����.mt{�w6���﾿s�}}{��{�d��Cź��͗9v�Ȅ\+�H���4eoe�Mv��k0a31tz|i�9��.�doP���}�B���hp��0�j	i1SK`{z�� +��*�gw�]����^ 	����p` �i�KiȺ��ޡN��Ъ�#�xKř�W����s�����/����z�o4�M"�����R�2�j8�<�An�qtN1��& 7݋QF?w�o<{���|mgqՎe��tqg]�ڦ���e	��$~��H����u����M��n!���Mx|o{e��O�:Gs����}��ޱn����4R��b����4� ���d�>�Pti^oX���������K�I��v ;X�����U������A�4�e�e�9p��K�z�B�<fݣ��X����B�-͡��v�wP���\!G�F6C& &�������o7���ף��N���~���,��>D��4Hnb����T��Щ��w�w4�oP���G���l��w�����n����]Z�ޡN��wn­���el�/��^�;r�W&Q
���4(��"���f��W(�趩!�l�nfs�|�"Q���]����1ipiUG�u�����E<�EiIu��[k""J��,�ե�����)�w�������Ե��$���À�M��G=�SK�|v���Y��v�:xӥ���D�`#��2��J�eԨ	եĵ��$�4vh�h1�2(%�`'�N���c�B�-͡UH�����w�U4�J��i��-��b�������c��xҤ{{�.�doP�}�{������	�wh�B���ک��}l����Y��v�6b8�a7	�0�4���v��eZ��P�KwhUW���wX����Ǜm�l�wsh��
�^ ���^��R�w7�]Z_E�����S�^�����د4�]�S7��t�ы��.9�n:��Ja�&� �w,�"-}�5{��r�X�7��1rE�K�9w��4QBI�!�Nh�KQ�-2Yt�f�f���fS:ƀ�+��Z<�4[���MB�(m�MVPP!���	�T5��]��0��t�Bg��&ͨ&`B�i�\�b���;	���cP�7Zb�n�.����;8d��4j�����DW�Hܔ�1]��)��jZ��]W	������B���׮�˫.�����?����dU���cj��5�;��wg-�����֔��
@��	�o/\�J���.���h��f\�-���2�E��4��6����$D�qA�Ŀ���*�ݡSH�ͯ��ul��
�^d���B-�)1wk�uW��;g������z�:[�B�>m�8@MD0ۂZLT�>ު�GshT��y��v��>4�woRbۄ�m;W�z��-���T��Щ�� �=�sK��6RP�pKp"b���Ъ����q�h��.�doP�K� ��J=	��k-�ļ����F5�Չ��z���Qw���vSBh��7(0pQ.	ln�=��
�F�j���������{�*�kZ� ��L?�Cf�%����_�÷�O�¦ɻ��M��K3R�oDq��\���驪��t*�F�eH6f��ƩC����[ݪ��`\@$����G�G�w����K�s7ZgZ[k�f�f�,���`I���u�
�F�hW��U���p�)�d�Meͣ��
�W�B���-�*�j��w�]Z�d��4!�Cp���}�}�b���4�&f{�q��.i/w80����a��]�xҥ��7��X�;�)���T� a��a�	�e�6���3�\b�ƥ �EuY[��3�+p�]�-&a��h"Sb��l��9yB���hp�}�xҥ��e#�a��;W�zD�ޡ3�d9���|�ى0�l�6&b��&c1<1 ��,�S�a��J�"��&�L�J�-;a��O})��v�W��YK*�u&& ��/f��E.��Fj���#���y�kmv��giM�����3��mz���"6ű�^mx]Gn�
��; �G�A�Ъ����x\�͙�G/(Tր����Y��j!7�0�4�����C�|7��Z���*�ݡSK� F��{�a�V����4uYI+�륎�(�wcl�ڵ���b1�!�&�B)��w�T���T�<>��*i����uio��"��!1J��Я| �g;�T��ꪤw6�w��V����
M�`�.�|e�9��.�}�=���v�}UIZ�4 �P�A�-&*k�>޻�G��T��m
��S~�B/��Y�מ��73N�M��{7PN8蜻Gu�Kw�%]��(�Y�'*�hy�_����(�SGpS�.�h�鮍�U��$N��kS��3�>�0@$�;�[�L��Q��m�Lh�β#mֶ�� J\|�_��!"
�-�V�WP�Ax 7z�ݣ��*io���ׇ�>>���6�MCJec6�n�ጻ9F,��k�iXsAm�r)��e�e�g�=>��v��2�nf���]���
�սp�����pKb��u{����쪍���T^�P��뵾\��&�L0!�t�wz�լ��)x}��ޱuH��
�W�8�"[!��Cn���wz��,����G^�s���7w�eZ�@Ǐ���
!���fm
�^ ��6�{�wV�oP����_���X{�f��R�H_s��uI��wd��9��qv.`�<��W��1z쑔��3�"�|8*�;�VA75��ϟ��>x%�(L��5ښ�A��4����l0��Yi/b��@+�ˬ-p؋B��6J��i���=��J����+!��ElԄ fk�qw��O�,v�Mvը�&X�6��cH���^�{&�Db1l(��:R�4�fn%#Sh�E��[��u6�1�,nV�25� ������v�u��L\!�k2��Vi�����,
pm!Ŵδ3�����&d�����	aB��=�x_q�l��ldv�j��J��pC��90�c0Zͭ)���0�b!8i�l���h��.Q�ͱuk#P��6�z�U-�1ȓXp�e�b4��z�������Y�뻱�K��	Y��FpKc��E�lw�)���}�{y�����g��0l��� ���]�79��+����	;�|#Dx&�UPo�\���#��
�W��.�1��I�x~�B���zŰФf�x��h�&�&�fl�
�lچ���g�3�Q��%ʨ��N�� 
�f�j�������p�nI�գ��(�A���W�c��CAHa�ɹ�BJ��j3lF@�:ʎ���kWe4&ʅ%D��"����J71<Λ��읠�F���?;����m����7h��ͥ��L�m�۬k6m�C;i��[Q� A$A~�<�}�.�=2�(��+��U�3Ϙ�AN"a1N��P��ov�x}����f\�	����D&�mC%'w|>>4��}B�.3dk����X���5q,&Jn�tf�c}�sk���Qy�B�.3}N�����d�NZ�9���k�a�eE�k�ꬶ����{1���_
��(0���aH����
t�6�U#{��V�7޻�^�:)�	4��CI��W��/���c��xӤ{�B���m
���{;\�y�����,�ػ�wު�[�w<#�Z+E�%GmyJ�J�;3y���R�uxp��Q;V�ح�ҫj�Ӄ$��D(Fa���<��T}��[��e޷�g?/N���5�c���Q��x{���YSbr�DN��<��j>�t�\�y�y^�	��x�q�\!�z�&a�G���� o�S=}LԀYJ3ۛ��K�e�/��]+{�7y7�"ɘ�Ѹɧ��zut�0���J�g<�n�X��"![]����Y�ק`��td�D�}��������N�Lp��;,lJ��yF�<�]����s^���;�8'�#����1}m���,h��*ܑuVO�`�"�]�7�êF�����<�J��J�����n����:��C�K�O��<Vǅ)Y�& ^\��_���$�rd����NC	B��b��[��&���{ ���z�ܾ=ǩ;�t9���m"{������ٸ�<6���v�ݜ�&޽Xs�]M�3���I�Gq?s�L�z����9����Kv~/�%���c$�E��g���'�r�.�k��2�[
��xѓ``
xoK�݀
Ƿi�Z|�wpC&����a6j5�3�0��E�@�}��zːadS�z�ڊ��E�I�O*A�娌�ч�^	�v�3�Gt�9m	����˸��C[�� ]�p�Y7c�>ǳ�ZX�h쉫��T��l�o�T�B�J�H;�^�ٮ��2G����킍;��L��;�{{a:/1���Nϛ�[L2����[}�6w���o�t����/��k"œ2���TN�"*���1�Iߍ9�e]�G�v�����H[�n����\9��J1Ꮦzv��5�h� ���$sca��6%3_�owf��]Q�9���<�=��'��=�pו%�3�bȞ���v>\��Xm :�xŜ8����AJ&e2kqHqA%�u�%[W4Z�5���j<A#�n���ׁvq�]�`��@ ^6);��o&�±E�G��ޠ"�(��\1w����ʋi1DAn!$�T�A�cS��$DG���V1C�.f��Vr2e��m��2y7Z#G-^�TJe J�a�ni�dmc�h^�ޏr6o�[�iɃ�wa��Vk�k�+�!��b|��٫���uE��5�zcype��
�so���?a}�a�F�۱M���Zo�s�[��A)��~#5T�~�4��9���2p�}�u���rS���ӄ��F��Α�6gT>>���p�k�F�$P�� �M����8 ���'�����۷U42(�G�A3���8|�(�M�݁�X���t�jCP�NNu�H����W`�wY�������t��qnT!��`���)�U�<uI	|p΅L^{���0���e�x~_�h@Ĕ��m�P%��b�(��"�SE��x�m
�[��.�sZ�'�L&Ke�b4�>_{�I���1W�U\��uT�� �KD2\Am�ͣ��*ix�������ƕ#ݴ*ix}ٿ3��V�4#9�p��MB8�Q\�ɨ8n*!���V��5�õ˩��ܳ��~|�B���ک�������g}ꩤ�����[Pp���[L��{��M,�u
t�v���]�ɎD��&�j!73��]�����U���]��5�#DA@E�S)BTw�������1W�U]#�S^��!��P�*�ڰ�� ��sa�e\�$N8���E^�ml��l�GC��<j��YoK�׷h��ȓ��������_(�df�t��fQm�˳kc6m��R�j�N��t�α��֊,����:���H�0و��4�7�]����Sƕ#��b���H�+��4Z�Ri� mt����Q��,�5��±��uXa��|��0��b�h�[C3�z�ioo]ݣ��< ���ޱwka�yy��,�P�*G��W��Z=���ڪ�3�Kw�@�� �ᨃ.��#������}���'�Fv��|�E2a4�LUx}���0o�\�j�������]F.��pa"�M�eBb�2;eO����b�7ޑ3�"f'Ч�)�ܦ����Ȭ��9q�e�]�[K�*���
�����5�Q�l��C����kh�s�͔p[��r��	;�N�Șˉ������Thn �'M�Aق��Y��s��1�ذ��.΋�-�m
F�(UD4�u�+e�,��[���f��^�U����sR�YIR!ĥ��ԕ�ڎ"C3&`�ԣ��l���OΥ�\ \S2���*�j�en��9t�YP�&�̦��1j���nT���+�k�U\���R��t��Dn�`�t�ڪ�	`a�b�q-5|��<�~w�
�+S�-;r
-�Zve�a�D@�Im�))H�<c��(�tr�ą���e-�R�L1����L̂:�� ,��8pJn��귿~��G;�TҼޱ���f>��T������!6Sd�N�գ�> 	�{�:���z�i^mW�����\0`��0�"LT���X��������s��eZ�zD�T�!kI"QpB�[w��o�w4��UT��Щ�����k�pE|�)��٥H�wX���t�R�2�U#}ꩥ�}������Qv��m�:;G\�­m�u�+Mc���-4�\�;B ���.Y���B������[O�
j�{�]��`ǌ4S�	4K.LU�Vv�~۹ddm�3�I��Ѧ=�"������R@�[�6g�/�"�ċ�Ϥ��67)��F��WB���.����\�"e�%G��H�؝dciն�ͯ��/��	���{vf`�d� ����e���$�dD7w||�e�9��.��ϤJj�(UR��י&l�I�Y0�Mp�뻤{z�M+������|��xڥ���PP&�Ciغ�y����̿���UM/n�U/ h4z� Dl�@��&6Ь1���#[�͝��T�����sJ͢P�0a��ͬ����]�xҤsw�{��^3�j���h�SB����W��Z���n����j�z�x|-n�G/4"?�i3J���X����%S��Y�׎Bz��;v�Wun^��8l�Wl�
0�n��)���(%`ʸ[v��X�$i���eNp���f{NF"��Cxx�QJ��i����;d�r��
#�@& 1	���H���ꪡ}陋�"lw�7��ww�>Q��1{����C�+�}�������hM8D�aLfgUW���S����oHs��7��daq�a vVh��lõ-v�@�W<�\2V#�B�L��W-.��Cf~~~o�w�O[�77�]Z�]C��mm>�
�KQ�0�ÂSp��������~��c>�X���ޱwk�O�m�x��PpSe"[NEխ���nm
�}���w]�.�w���w0i���l�,�����}��;��2׼�ƕ#��b��xת j�V,�?p�s�V@N�&{3��W#�R�N�A�]�V�^��e8����"�"�(�>��9�:{��uYy��1E�OGN@q��i� ���1��j�m�ΛY�޽��J���KС�D�Il]�9�U1����{3 ��N&�*�� �z�B�ZA�!��g���P ���CFV�1;R@�v���A��-����+G}ޱuk5u
T�6�� ]�9�U4����P*`�È)���{dO���y�*�ll�ӤG��W�­�S&8�-�	0ZI�J�oP��ov�{���&��H�+^f�!C� �$�w�|���n���
�W�hR����.�k��L�@M�,�n���{��׾ G��:Y�B��FO�:X<�r{т��\�]377K�̔�Z�\hL�4;���U�P�{DQ&nJ��[��J��{Z��gC�tb���ھst����U�=\��a����N	N�q���Tc�d7[�-J�Y��Fk]���T�0��k	�;�tʖ���%k��F���Q,f�"�L`f�([���5uó�I���
�heŚ�cG:]!i��.(�%�,q3M�#/���X��˸��^p�޴�j-0�RV7�5���c��]e�l���Ĺj,ѳ@���"�Z�V���f��Z�-�c���5нN��B�l�{�/��:X+fz���*� ��2��5��la�.qf�8,F��d(��EAK𹵾_�R���*�ݯ�|.��o�w6�����C�0��fm
�����Ɲ/oP��q�C���Kw�� ��I��m]��zfco���>�HN2�z��Tj\وp�(���~|�z��,���nm
��3��in������$����.W��nm���ܧƕ+ݡUK��xM�h8�	�$�,578֪�T0U�vu�3�V��ͅܫ��f��1n�oP��ov�i�u��^3�.U��M���6ႛ7v�T����e�g�~�vTO����k�y88c�ͣt�
�J<ci*�ڛ�d�d�X4b�k�aF��E�.4B�/8X
'
��On(�β���9�f=��T���P�KshW�]���'��m�ZN��{޻�G�D������.���+/@�(4Se"RV.o�Wzź]�B���ک���{���^�84�H��C�DCLT����wk�}�xҤov�T\g�)�g���DAB��m_T�2��Xĕprh:�-��� �,ɜ.1LVId�y�7ޙ��;�#� &����w�8%�&Kd�_�S2��;�_���z����T���pU��@(�%H�Á	eͣ��
�]�\n垊��Z�,��7rq�8�:�*�%�=��t7�T0N)�-P�I�ZauC��ѽCn/�2�S��3�fe��/\gQNb��f��#N�8��ܛ}B��+cwl\�ΖJ\Z@�\$�f��|�z��#��SKwj����ޱsK��Ɉ�	� �[$�f����eK���Y݃'G�J���*�w�v<�
�`y#��Y��aX�&�Bi��Մ�h��F2��5ٓ�K���q�n��wUU#��*i{6���1��|iR��x@�_ͷ(N�ͣ�"}��	���*�g�fcwfx )flP�Pb�N&Ø�oz������}�q��!���)��N
j���;�UM�GshT�s�j 1����\���|�
���N�����u��r%MA��AAXm� áo��n�+�c����!���S|�i�_�yo�ϻ�i����A�P�:j�Ezס�B��B�
%&iR���6���Z�X�j�hUR7�\ �
�BSCm�DI��Z˴�p�v.1i�t&���r�; ��"((M!�V#��
�W��.�o)���a��z�ե�p<�0&�()ҥ��+�|�9�u4�{޻�G;�W��U����`�M�d��ݮ�T�����}��z����T���U��i�Q'S]��{�̸;�Hs��w~���S�J=�`w�L�M��m;V�7�S�Ǉ���F�}2����Z���������?� ��uuwkW���A�y��q�p>�����]��;w����:f�"� ����  H�2
��H�2
)  H�H��`"��# � )"�(H*������ �� "(H*"��ęE ��"��"�	�" &"����� TAS�@9�̢ �"��� �*H(���*�(*�b(�������p"�b
H(����#�(���" j
� �"
��"�� d�"d� j� .H���  �����`����9�"�F���`�=�� v?�~�*Ȋ(H ���ك�?���y����������!���������/���������d?Y��=�_?��h~������������_�?��z�ߜ'��?�����0�����@�/��x����9��O�w��P���E��f�G������������h���������_������_�O�)���TX'���$K�!��.�� ���4�1�����d0`���c	�D����n��'�L�����_���UE(��"� �H@��H!�1 �F�X�D"��$B(�b��$B(�H�Ab	 "��0BDX�@R*��Db�H� �@B***�E���D��HD��"���*H�E�DX�@H�@H�@HEH�b,  ��D ��A�D�E�E�E��F*"�*�A��* @"	�$R ��A � )��(EHD	 )�E(�E�$TH�@�$@X�A�$@X"@P��
@V(�P�$E"��@(�A�$@�A �$D"A�$@ D�$H�A�$X�A���D@"�V(�Q"E "��$ B(�PH�@@b!A��(� �E�A �P��X�@P�$U"��DB(�
B(�B(�B"B
X	�$(�R(�X�DH
AH�@�AHA�DHA�@�AH�A�D�E�A(��$P ) "@V�"@",QH�@A��(E�R
P�"� "� ��A�AH�EH*��B��",U�$@"�` ��E*T�$Ub	  �A �B(�D"�(�b�(�Q�AE"	�EF X#U��T�$E@�$�H�A"�V(�"�"@B��$�$"��$�$�$(�B(�B��X
E"	"� � ��� �1B�P�� ��E��� )�DR��$Pb� �AR(�A�$b�(�T"��@b� R @b�(�Ub��$D�Tb�(�D"��DB(�
�X�@�E`� ��$T�$(�(�X�D )"��$(�X�DE� �X�  �@  �� !��*HD`) `,X@HX�e*�:�N�K���R�R�N�J��R�NR�N���+�}�u�t�Jw)�\�)�)JJN���*)(�*r���t��������N))Ҕ�)ʒ�������(� �R@aY E�o�.�����1L
�Y�?�7o�����PPA~�A`���������������O��?k��G���<���_��#��?�y�o�� �"�����������?���?�?t h?@�������A�d2'�Ӣ�?���!��zh?�4�y���'��+�?�����\bO���������~���?�_�N�B��AUD�'�(( ���'�#������s�d6�����xw���_�:O��`QA����cj� � �0�/������g嗹p�����6��
��A����iAA���(��������栠������?��P�Q\E�!�ca�t?���Xc����?���~/���1�c�	�L�'����( ��?�0�����ࠠ��c������~�:������m��D�<�� L&I�d����?��Q���?��"VD��1���9q;������/z�c?g�~,�s������x? )��������nG�g��C���C�������p?��4AZ�����������:L �s��.����#X]�C����p���80_�<|��rE8P�"Bx