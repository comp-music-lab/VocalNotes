BZh91AY&SY���~0�߀py����������aG�Y��!�   �    h       
      @ �(     (   � 
� @�z@*���(�
R�P
P��� @�PE���   �I�ݥv�>��Ѷ�!�n�����vt;�׻{`��p�:�@�J �me���5{�޽���U��C�8m�P9��A� nÐw59��`�IT*���   r@\<\Z��f���wb�3p+�efhMm�{�]�J�x^��{����)l ��]�0m�P��`=p(��Ѡk{ z���   �H��{�#F�m��@@k�H�݇NA�����4t7a�
*��-��r���p�=C�{i�뽁�;n
>G!N�=wj�����  !wP 8^xm��v��q��ZϽ�zk��z4빨`>�PѻQ�AIJEhoq�^�]�ltwa�]�"�}��7�����T��p   e]����W�׽�@-�ZX�[<��>���=��w��z�A�*v�u-�]��[�ڏ-�v�=�r���ݽ�p^����2m�듮�  P  � @�  ��   ��*U#L�	�bL �� )�0��J�0 #L � `�0��UJjm%  0   10f�
j�P��b`�M210 �'�RB��� � 4    !j�bd�B4�=�����h�P��&OT�/������_ٽ��[{.�"������U@�E�*��D�"�*�h���_�O����?݈�0UN�T�o�*��?��@C�w?���@ܢ/q��O������?@��I_�t~�����s_���u���3� ��z�v��k��g�;�|	���yu�y��Sw�Y��v� 	;��Ԉ��'gm&��p��#Z����8']m�R�2� ��0�����d��Η��R�i��[�d�挓�_v9+���WPb�m
��ig.�r$n�L��2���>��%A*	PI�	P³����^;��q��Q��&����,�X�X�&���'pK�(�UWU�k�]��q����l2��wf�:��}G��}��f(����n	�>Ͼ��ϋ���R����yދ;3������� ��x��l��������?�?&C��Xh�C�Q����|����� ��<l��F��·�;4Q!���k(>@�Z3��r���6Sr�q+��c������l�٥�d�t�'M�G��g�q~3v�1�-���c�h�w�F�[^��o��uU��棲�\H��m���Oz�|�L3h���{^D̵�f��>ja�2h��p(����~�/]\�m�H�p"��ƶv�[����f|�e�P�Q����j�;4h]��L,�����O��[n��>��{V���5���rި;N2�b�X��j��%i�����Moy+���w;�9��8Iw)v�;L���qlͅn
���e���y�Y�ɋA2�b�AN�x�8:s�#��l9zsgᣟ`�?m;`N����MtSo����H�q����R�$]ҠC�{Q�x܏�H$����2��u&-��ӝ�ݳ�0g	woK/�fޮ��fӛ���V���֜dgM+dۣ^�u]������RW^k�&j1t�tc�Ю䯁G���`������|��wU�9���l�6�lW��
,y��ׅ�;���� tgf���gwL�%��q���k3w	���� qIo$���ߝ�3M��vl|r��d�������c��cq��0kص�X��fh��b�6�}�>J�[Gz.�Ou�\`L\�4��v��)���c���9^7����OjN���N��v��ڰ�m�lX;��"�a�x(��x96����ۯ�b�M�t���l��@�y݉�KJ�c*�ٻ齃{�8��qv-��.;SԟF/l��x���6#ˡ���r\V��;t��X��ȑ�*Z��S;tA�.���+�$Fݳ,�f���q�@x �n��l�f��08@�t^}���_����H�^SbP���w�ܻ1Q�����y��6���T@c���V�wmI}��b��=��n�c˛��:j�K^j'V���.�&���W'�W0��{s��Lɪ-�F�H�i���w8�yRŹ�oM��9����歲�0���ֽ�N�<,yٷ�Z��QG�m�7�c�J�x�|;UPȒ7��M`�-�9)W\�E�E��-�oc��`�.�,����&^�����hE̛׹���Y��@�tQ�|-<���	bG�j�!f�c��p+�Y;S:���0�q����)��S��9М)�v\jn��}_O*�	l�R�u�wFL]�s�y�ͤN����!F��sSt���᯲�i=�=��-m������sN.���p<��?X�)�
�*ӎ��z��b�nkYT�ó�ԤgKu�h��$R9t����/�����C�Op��{�Y�Gs�O�A�vr��CK9�FF��Q2 FLqw��\w�W���z]�솔I�� ݻ�f��q���(�:��X!W���3���ew,�wCΆ��Ү��x�g����0�q��ƨ�V�˯:��m�"֓�2��;U�+�{���.��R�{/r�ƬU�0�{�w�9�b�'7��yv�9���4r<8j b��=#��{����]�hkf�q��x;Di�!a�[�n���E]{&z��c8oop���v$Hgu�{�:D�z�Ҁ��ߞGBq]f���!�i6���v{��,k�uk�ɲ��q�'S;';"���Y\�������^i�������p�v��;��Nj�h�W� �e�N�ގ���&K�]������t��2�ޓB���2ےܑ7(8�M�R$�)��{��fǏ�(93£���2-����w /qv�cw*�X[����*��k��1�����
�[qϤ{��j�l�p�=Gp�S�q9�ӖK�����,T1Y�n���j�u	{r���u��t�v� іkl�%���Wi&��da�����x�d�&ssv�N�îQ�un>�H��y�c5��ҁ�;Wb�v�lY����</*���l���Ԟ#��z��&��͌~��1o��#� A���4Pd��=Wqd����v�S���=���a�3PՆ���.f���viU	���dv	��Yn<�r7Q�dƬ�m�sw��a�9��O�����*�ݻ�vR�e'�B�~�@��x����y�0 3�˚Z��wW6A����h1V�3r[���J�o����=]��}��lk4ep&��'L���P�$���1��@��o��ϻ���7N�����L��tlP��Qb�aɼs���ZP�#![��a�w,��N*�^>	� >��ҥ��5,۷#m�d9��O=���hHS�L�{~"�s�������iڂ;�^ı�{o�, o��{�,�8䇊#�m���=�&����,})��|s��iI݁��a�aOWi���J�Dj]X��n�����-\V���X�kK�뇻u�F�{'U��$S� X��1a�T.��3�M��6�-����-��(��@x�x���͜�f�Ц��{5\պ���b���_R�s�l��X��0e��7��{4pӜ���`%;�9vώ��!+������u=a�	��2����syti�R�!��8�M��&G0ՀQ�Q�t���c~�ٻ�а�P�lNi=��Z�ѹN�zc�.��,���p�"yN/o<��-�S�^���9\4��Oj�L&��'ol�8�t��9d��F*��=��!�^u�qY���������k�Ch�z#���tzDD�{F9ynEz�ћ�����o�ʹ�4�Ӄ�RH�C�Q�{���BS�ȩã4U�ʉ�8^uǮid��d�v����$�d�	�[�u�ӺтTv��Gp�Uu�V�S�F�!�wo]=F����ߌ%���K:i=�uokY�z��7nn����f�5m�x��!�66��&\����$�W�h0��2d'n���˞��9��E��$���ʫu��@��wRMz1杜!�6�U�(.�#���f��� _-3���U,���7�ʭxx��x.����zU.��u�<�X��\wl�n�m�4հ���x�
�#�
Ŭ3�]�nwf؆w��K�vA� ���
�2u�ڰ�s�$&kI�ӥ��`���At�S�	W�)�j�F:a���ݝ+s��ÏE-jG*ݼ�<%h�]�'*x����1f��atSP�k`�.]��`���7b�� 8�-ͳ�����.N�b���m���w��9�Y�V�"�F�� :B�Ï�y./����6�H��4�whP�T\=;�mi1v��!�%�1�V���=w�؝jܭGy���Ӈ9t���_��]JK��g@���v��XN�����^KqvѴ �s6�흼nXp��[�	ق,k��P�9��ӧ@>ס׬gs�� �N����
�7^˝4�V��q��3�I���H6@��K�ҽ�8���.88�N4��H���p����lɽ&�7�xf:8���#V�y���k�R�d��
�(#�=R4��;MYU�ƻ�v.)\��˽x�wgnD!cM����$�ɭ���ݠf�5��:f��Q$����d2
{��i���_^�f��q=yQ����{�<;���0�f�:��W��>k�I'Mː�l��������&��V��^W�u�Z���>�5�w��X|Myr���L�Л3�Qr���ii�D֦:r�r>h`�^@���Ҵu��oV��ޫ���E��庵�8�>��z���87��K�� }yYa�l<���S*9�Ƿo-��[뗞��0t��p}�n-ʻ��vi�#�w��;e�o����>��ɓ_	qr]`j�dOg-�HwG|�eY�k}V����wv�g�H�$��w����<Mb[ɝ �Ŷ\/d(Si���7S�$��Ɛ���P��;�N�gU�4-թ�Ѡ��ٜiq�V{,XspgGF�l<0z::(�Y�l��<,�G�d4gR:�YetPl����٣?�n��������~�~'��}>X�;=�����g���]��@��ދ5��/�n�u�n�����j4݊��X.��d�K��,���h.zǞ�{\v۩8k���i����M��C�W8y��7&�����e����6y3�Ÿ9�b}����Q���O	9�<s�݊�9��l���<3��Χo6�u�=�n�+��\�.�n��!Nnz�8�Uڈ��Gb��5�f64��s�z����Q�t<�v#��\6J�������t�[��(&�l�Ík�幺P��/�hƧ1=�.6��zw&��:w=eP�q�Ӎs^ۈp�U�6���� �\>�����ԓ;�rZ���zn�M�w;�.�f��l���4����L��U2�R����qnK���X�#k]]���!�n�sϧ6;���1`�v\D6d�:���ζ ����r�3� �w*j񎻮����M&�<U�zݰv�s��nlg��f9�o6ۀ�3�óYS&��g�4�Ĵ�.L/>8�';jx��kpa����N=�����t\ ��v�q׷n�:�cgR�a���.���w�=�vs�wh̸{2����r��^��]���9��k��kc99\�m���W��Z2�ʹ5�hq��7Q�@�L,��A��b�^�z��|wZ�|�N+������D��]�� ��l������k{��ms�u���R�<vJĕ�pm��m�1�caJy�R��8n��x\�x9�M'ǭSu�ls\/6�r�7K�<�ܭ~PZZZLbj6�kv�%��O<8�dq�z���*���vP���Mk�Y�ӫ+Ѯ����^o8�rv���mC���=d	wE��v�����dM��W\.�\����0�P�������$M-TԈ{����}_ ��o��r�,?���C��Y��[+�8������u�ʴs�͍vb��1�͗X��^܎'r �H��m�c����\cY��ӵ�ٸ去]m�l���\�E��Ӹ������^n�\�� ����N+6L��9����Sm�60�F�NẈ��`펲n,N�1��r×�������Gb{�S;�����cK�]�{cv�7$�8��`m�d6۫�n9ְMمݰl훍۵��v���W����D�y`͹���}�7ϖ/OW���:9;�����vϞ�n�/�<lܹ����;�.Z���h��v�P��sT��
��k��6Cld�:��u�)�^%�ֱ� �Z�r���9�[|O��^����#�W��^�r�끹���U��q����V�m���΍���>�sݼ���w�a� ��n�A�X0Y��9kv�բ.��7(n�6�N���Ķ ���]I��Y���9��vxu��9]ض���
�s&�=o�����j�eݝ���u�M���S9�F�W�2�k��eX;n#�^���u�i�s�r�͓�[Q���$벛�W�gREG�͘7U`�[�e=NA���(���ӷ�)S.��\%��j��8��G8ޞ��]�K�ՙ����ۗ]F���e��#�kv�rm�Z:x���k��v�mvܴ��ۃr��C��\�q�\�����+�8��X�М�&ծW�����$*ԏ�n�i�M@�l���ܤ\>pX�ì�E#=��ɫ{�k���w��%cn�/[�n����v�Ʉ9^��c�<6�om</i=Һ����Q�9�\���k�[÷O\=q۟[�����v��C7G[��#�.^{j��2�N��s�v�mX��Ѭ<\ay��������[�{o#ѷP$q�<�;��v����d7<A׆.��x�����q�F!T�Mq�zl�Ý6�u���{M��­�4:�uۛj�gq�n�O<�wnL/6�jvq��-G��$�q�s���1���;�\��t=�|�y=�6�. ���	��Ժ-��ߋ�8���[��q�n�xy��[�M�xy�'�:�:�����i�@�[q�j��,ݵ◣*�s���ٛ���J�p���5��ݢ���squ�K8��d훷X��G.N��{s��g]�;�=�67նwT7�y���Ԙ��	:�Ry8kPu����BRD��W����8��U��L��m�u����R�K���L`��s�=��2���d��`�bo'����^�R.��mn�s���#�{Go5��IĖ����ϴ���q�SՐ9zn�ac��������9W=���n޻Epٛe�����C�gp��e�ƻ1�I��W�Tp<u�pkc��v��q�\Y�;�&Mru�H���-"�D��B��v�ls*����v}��Ē�;m:b���?;��gqWb���*��lr-������H�ji��mnʏDy�uMr������ �)��5Tk9����[F]��c�����ۭ+� Yb�E��޹<⻆J����s&4��f�t\o�7]��>6�7F�8�۱l<l�_9۶���՟j��펺7GG'�r\8�z�� ƻ8�^q�Q��A�i�̝N���ჴ���wdw+��d���n��1�/`ɻ�W%۶��:`�5��l����H�m�Vx�cv�1��=�=��à�˳2;!v��j��oX�Ǜ�/X�m���:�c��ݮ�3s��wM�s��0Z�;��3�l3�Ӯηr�N�f.ֶ�ѹ�M�óⓖ"wt:�S��ݺ皉@�9�77\n,��=C\M���|������ós�ǧ�hꝸ�<���~b쓕�&-ۨR���ݧI���B*%�ʤ{1�Є�v�2훷���m.�3�4{E�K�� �=�1rP�ф۳p��zIv�Xx��,���$�p��n:������.�:�/^yd�}]���8K;lY`	wb���-s�}�mu�����>#�rܰ<�m��:�~�I�����go�u}w��}�|[�%���r�]\fի��w9��u��<E�\=rBķ��$�=J+����Z�;b�F��}�ѫ������@Cw�:�y�D�WT������|/���s�ԗ���2�U��&u�_�)� aٳμ��y�!�,;U8W-�w��-Şv��S~]9�wun��H�܏�j8E�ѻ����:�=��A
(�B��Μ��[}��M�<�oO��|_��\>v!�������/����HnL~f�v_v��h �O<�~<��s8�3�����Y��ȼ�#���d��{��=o���q�:R��ゼWMZ�5���Y�9J4� 9�<��]���~(���ݒ�p'�N�Yj/=�|<���4��"�U�z�2��[	b�e=s8b$)�ůb�+�`C�1�ș��\����͟�DԆ{�;%���q��/��h`��gӷ��C�5�r�3��Xnj�f���3�P����'e׸6o?��;�[7$�'ݜ]�{+�k7�V@%������E������x���v��ս\\��.�۱�Y��e�� ^z][�>H�٥I�!���0�+�y�5���]pa�����N��Y������Fj��d;}t�L���m9`�����vE�fᓕYz5NJ�ʧ�"3a�5̓�o��t����򛩶�v��֭�^ ]�+��kc�۞3�B�C�p�����x�ŉo�+}�̈�u��ʗ��Z)�,5măO%��}�oۨ[��'��=sq���UQ��G��u�(nH�h�����`{����=@�`�>��釽��Mݫ���� �$��@���L̘G��6k�[0�\�r?4�w��ֈz��	��[��w�;B>��6���~J�y���sV�[��w�-T?x��7�qkw��a��f���a�U뜾��������ܔ2u����Ž���n���G�� �<H�)��b�9�.�V����Ǘn���0{�.���r���!�|-��W�n����!nv���3�6 �>X�4�EŻ����h&Lv>:��u�=��k^��XO���?-^��!=��x<4��=�׀�F-�����[������[xz�8n��sq�FVL��SҢ�d�}q�y{'�=2�V��qga�i���'����>>A����^�ݎzc���^z���5 �K-HA������ ��sh����p������Vn��!n������<9���>\ה���_mX�u3��Tj�Z�m!�dJ�[��Hۍw�wH�{�"^[O��ݙ=�/S�]�X�7zzq�W�Aۂ�90��X\�ȉy�����V�"�sql��x7|N�&��n}M�����Y4��,���f�Ek�{=��31��τo;�כ��f��UeCV�(=��y5��Ħ��m��n���M���x��=�<.r=l_r^���ʌ�4Ι0"�8��t^O	��y<�3^�z��茒����FC�Myhc��;�&�徜��z�1�E_�M,�F�`�nѹ�����Q?���<J̳�ȇ�����H(9���� A��8x��k��;N���Q�_��,�;ȣTh}D	.=���bQ�q���"X�G`c^(�cFVi��15�10�У��7j���	���N�J(m�D��e�A���6�#�]U�v���<��[��+�s�w���j\w��$�xs�.[S���=9'=�X�N�}�vv�r+=�*\F����٪�<��n^���t�5=$gx��(�>Ƕt�{U:�qYn�X�B-�W����HR�s���(7}���1���£�b��3ʝ�iY�U�d���%B���ܠOy���#4���e^���P���5�,�d���#NO{������m��+�3��`�o�vq�̈ٸl�'¦.�&�2�4���Ո���Ft�q�il���獇
�b뽝}c�X��U�<E�Sg�7O��Ck������1s�Flg�ś(�{_=���u��ry����Q�9�ɹ���̻�Z#t�Ϧt�y���t��wb��xꖪ�+3��ǠLZ={�H��u��
�q�ˉW`�9a�n8�;��v����~c��ae�(ɾ���^�����;&@�Es����w)7y�y�<Qo}�XX�f�/+�ƹ|�)�eP��R���G��}Ew�ڧ8�>v��u}�!�s��.����0=�T�8�T]�}����|w���j�aC���W][*>'�k�bO.7��gT>ݰࣼ�hjr��B�C�̶���F�omS˭��oz͗;�t����<�@G���ޝJ؜��_��op�;��؎i��aCՙ��t��y0���t��ӽ<�:�B{=dTM��/k�/p��V�s��=�,��l��<wz���2���y��{�bF��6-Օ��=����
�ww�g�{ײs[�%�͞�|����yKS�:������c1Z3^Vb�W�P)׉q�75����:(�]j5�G.M�qwxA���yj����� fߎ��ޤ%�Ш��']=:IO��V
�WY��Ց2�T2����F��h-����!�$9��#A�9LD���&�E^һ���j��d�}ɯ�g;.u#�M�a-������E@-�͗H��w;dVb��$'�X����z��2u�D���3MxT��ma�fM9� ��V�t>rw�#����ޗ��G,6�w�L�����v��cp�wgQ{��
���;;�G�$�><nm��г�r��iy;���7�A#�z%�c��v��
PDa��u^Q����7!>H�����;�;�($�3O{�i�"�Ό�����/2{���u�{ɑ� �W{hRK9A553��n���õ���?��
�sC:ȟ���}�o��+J�E|q[�"�{�%����Ӝ/Hޗ�}�t�m��7��F{|s����?J�͝t�x`�G�K̡Z-�:��-���f��=�M1^�c9F�>��_��IŔ\~Vt�ӱl9�L;�5�<��	DmnҵG6{r���<!�#�0�<~E5s����Ovl���<�z��'��w���\-��>���\s���}ۋ�&n���ic���OpkN�CW��w�x�+�)��	���J˥�y3�Mhڪ��.�{ݜ�_ų���,�}�w�'i����X��W���g�;1���'�����}->�����}�>���5�̫��F�n>�k�c� <=�q:�~�y�8�|q�=�+{�����Pԥ�Ho��=�T��'{���S�F�ƞ�����~�e�L���	����6 �{k�aG�7�/�c�Ys�P���{�q<���1�{��:�s��NWϻ����p�6;���y�2e��+[�Ǡ��)�� �܊���E;^v�&��Ó�7@�\��׻������gV����y_3��wIF��̧� ��O	��wl��{��ޣ�p}�}�Q�w����~ߴ�r�Y��$\)��]�7�I=�{����P�j4�z-T��w8`���+`��o�{67�{��4�lɼ�E�x�E���V���Rs�"�m�6N<���n�Ѹ�-u���v���H篙�/`�O��^�)e���즹��u�R����wD׵��v�]=���^�z��S�/7��{�L���:�F��j��|�mİ{ Z�ϋ��pXO���NP���j�Jy���L⹿B���K<)nOw�����m٩ۓ���������Hl�l�ʸ9 ��f���P�����z�0���,��˫����A��wX���Y�o�㰃���\D��{�8�Yf-y��[}�pl�n��,x9�o��%	 Ncdj�	���R]O�e�K�7�v����b��/w��h�p|�^��ܬ�=�_3~��z�L�����w}{��^�v^�]�yJ�mBq��Kvr[�D����O&␆�P�&]�dcz�-���[�����g����D���K��B^^�M�Gwd��P5��Od���cUS�C��j�<i�;�����kڔ(%�*b���]n�򞋖^A{5QI܍����jo�v�v'�s��}�f�Vz VU�$;�ө^�����>pG.t��ݯ=�n0a���V1�]�Wb��^��<v��}���',u��x7F�/6��٠�7wۢ���}�u';���]�+��|��{ �r5	$xn7l̅���i�هr��4���<�%gE���'��nV�ެ�C�w�U����9�lc�ܽK�C�Ž�գ̞�{x�M�^������}�Vv{�R��c����p�Yf����q�z{}u[SI	�%�Ȥ��DP�K����E�Qܲu(�j!�w+�SF��>*��3�r�h��>���y7"{7ֶ������쟷�/�|�T�I���?�?L��G`p��t�>�YEC ���VG���欗���4�]�̼��݀uų��n��:��g��nz@�"��ۮڵ�����s=��v���z��<�n�8lh�K����\Vѹ稊�۟3\�e��C�q�b�뙧y���\t��'����h;����[nX��������ۭ��:�a���n{i���G�)K��]�2d��e}�����t�Fysڸ]ص�3Ǘ:�h὎����ZCp(��gZX���+�	�]ݽ݆�㹱g���Llu����]&�d��R+�7e0��Xv��n��h�s���v�=��/]�^�<)	�D蜷�)$��v�m%ɷ�]��D�����[cݻd�%^�؏\[l���9��w.v�+��YN���8`��v��z�n۬��mX�n��vm۳���"m�� �%�0&��dy׵P�F݄ �>�q Ǯ�NNwvjӱ�v�Z�m���:}����M�;�.Wa�ɎxkM�۴�n{����ג�n�..-.wn	�x�-��u�v�6�W5��ñ�k�H]�Gp�ٮ��:y��x���G8�"ݨ���7���&ݺZ���Y��������1_�����&6��v#�6E�㪩���|�W��-����3t�]�ð�{��@|*x����o��x�}:�5��U��j-5�F��;����MIȣ�t���ͣ[�>���G�g"ħi�s��8F ��v���ͱ����"���&�۽��oyV��9"Z@�Ek�V����뫎�̏�c�9����˕ƜQ�=H4��W�t��)e*�}�7P�%-%[��'snT���T`�7�Ơ���iҫֶi���@��Ҽ�˹k��S�u.�]�ӯu���J	n:�g0rt���d�N�b�K�gU���[����:�g�SiiβK�ϰlN$t�#�@�!/�K.�;���9�֚��IJMB�Q�6�;�T�\j&� �o���h��?8ô��� �	�a�-�C�	w� 1�Q��	�����Tν\X�]I���i�NyY%�Qg��{v��V�&�4�Ń՝��u��C����:]�{n{E�g[g�]ke%mk����k��W;��rO<s��qWm�Lkq��u��*��lZ����u�ũ�q���w<���|�^7+�U�@Aci�f��Z��8��dL��j
0C hQ����_x���3,��H?V��@�����b��OK5|��q�#����Fv�D}
$����D};��v(,eY*t�D"٭��{����7�
  ��gp��H�I2��7��ykOs�z߭�Ƹ�� ����X��:v�X���h���W
�����ɫL�>��AN�gxn���D(fM.;˵ÿ�gq�ܟ�c��Xb����f��z�%m3Xud�p�l����Lv�ܜv�h��$J@i Df6�nLJ��J����7�~ڶ���[y��z,ɥ����} DEPv�I�l®Q��t&�c	�	ˮx`��S���:����0a�L�A�	gn����6
�<��cT��B�6��ߦ�������ڡXVkPa&W�y� ����Vfog�����--G���ғ�u`�5"-|H�!F�ȝB#���6��Gb�:���D�8�FD}�f h}"��Deu��8P�$�6�X��d@�~D��G�@�B�}�D�f�W��#�ߴf��˅�nb�:��LWE�9�E�Z�l��~�n13y�y!����D�O�(l�ȞנW���HbK[�K�}�8	ډR��r�B+,(��'k��ڜl7��Z[������(N��-�glw�e�s�r�� ց�@���:C�Ͼ[ϻ	�]�!(�Q�Y�1�T,6 0$q��������O:6�h��+6�v�]t��owDyo�D�������s��~�M�\��" ������2���BNr���}��t�s��I��~C�&�Tr V0�U�P�@0��n�l�F�M߷��~�R�gV�!]lF�+8�b�*N[{��*��sy��B�8�6�p �
I�L��g���Pn�;5b��S����7ʩE����c��"@0TN�g�I<t{ۚ�s��_^�X�#�JS=�9�ۡ�*��CT�-�{�l��߄�ެ���L����,s^Pu���*��VGA��Q�d �P<[����ہ�q׎5��n(�[�"��U��ۓ��i81���suYζizz��Kmw&����{�R�����m$W;V{�[i����(��ee�pYC"Ȍ�H#p����X�ra�!r���%C��s�^�_F�.�=�a|���PL�f��8�0]�&j�&�O�"ԓ|��!^0���T��
��S�A��JN�Df&tuMb�]a�XZ���&�z#ڂgS����+�G�� �'-��X��0��BB���12:u�ܲ<���[[t/#m
�bQB�,m��}���~�8Ю�:�N�(6��90�r�(w{�Q���[�1W.��}�@ꨮ�˱gz/�f��!������ x`� j#s�Fd!cnWR�g�"*��q��{�5-��%Z��a��H+GD����}�uI5�������P�/ J"I9���f@���U86>d�Im�A2�h��{9��1���jdV�~��y�=��%c�c&�_Be�i�'y�B˷֦jw�gM��i�����7�U�4�P�΄�׋��2<��~��zE�oq �:���Y�|�Y�*�Vmv̈��vr���(H�J��u �kV^j�y�W�]���k��N~���o��~��n������pZJOs��F����Φt~�����'Q����8y���=F MT�(�Z�r���=�����J�a����l�r�f8߾	V�n�#�=��5�(>�)6�T�$oď��Y���^�:�H4������LԷwHq��Q��={U�'8А{:����+�`9���y[�Ȯ����� �F@�dn�Uߵ����=�u+"���Yn%��V�X��!i�`7�D�6��>K�5%q�#:��W�vXF	@��AٮJ�~?fc�͑��&:&n~?�V�+������$/�D�Q-�=�:���]�&�2D�<M��N�wD���)��]��D�G�1��pw�b�u����g��`��5�D��dQN�]�:n��;c�Z�=&��c��;��E�{s���;|!>6S�t����k��9�e��A�t�ѭ�`�m�+�{;�u�O=��Lャ�ϨؙZ�ל�m���m�\7��K���D2��m�:��di�;v4M�e����u4���e4nC����h����Uz�8;=���!Z�6��u�MY�bU[Z��Iv�>�Wވ�����U(9zR�$3	����}���9m�SO�	F�gBe�e�g��2��J����\�<l��[l�C����nD5�./~�sgz۶Y. ��I5�������`��iy7����ݴ;�+r��)sM�P뇃0ٍ-����\�V�d|)���۾HC��Q7���5�EuBA�e}K-�,��:v�T.�1�8��.�'$G.�d��&��וf�њ�I$£Q*���$:����V��@���'/��g���7���ͳl$_�)��r��K�ΩI�xT-Pa!	I�� ͉7m�S�}�g��
�Im����ӡ�s�	!�n��ӺB�
�B~&=���"�%>�E�ۓv��>T�\\s�>��
��v$7t�`^:�}�X����7w܇��iU�J��P
�<zz�˽����3��(X� >Y�i����&�y021���*�֦�d��m�qY(1�zd�x*-��P��$C¦v%�v�^��]�<���K�K��ȷTB�W�M�E�`�W>�w���}�G�@���{D�������܊j�9��2*�w����4��h�?�E9y��2�$9�lˇ��ym�pu�D���6̝ywY�je-Tw��rf��Î>�^QҔ>�6�^����d6�n�	;��ղWʅ�������%\���=�x�?���@�e�����-���t3��^GU���[%�^r_��Lth�1[$jhE��Βj�w��O����{·�%�ĭ��o�-�!7uꋏ~o�<i��F'���="���?-t��KPg@��1�F(Z'AUa�����I��Ȥ8ՈOx��*��󉡄���ڬϣ6�L��k'5P���-=blʭͺ�XD�	ŋ�>w0��A���pC@�dq�\Ѻ
�/���Xw�5B��lсuk02��;�l�l�WUY:�w.�Ҿc)l�WR�D�q�l��k��QG�y�
�^�v���Hc��f���C�#� ��FkqQ`�2���-��ISB�T��!۸[�pIـ�o)l�r�	��w��9x�q�G���iZ��-k~�����oJ���&l��y^i�@'���5�<7� }�h�d�o\�����V�F1%�5f��C�4"��{����,��$j t�i���+Y�l���\�c6�]���t׺p⩴�:s�ei7�V����@��	|�/���G9:F �*�ݙ4��I#s�o�mp�Z:���Zd�CrG���f�!�BC#o�����.hߵ��kΎ-��#�sB��$<"�j�B$S�5N�
H �y|*#Dd�0.�<���W�[�G�����*K���;�C��cQȳ����/�x���ƃ����޷�t!�N��9������h*=�O+ �j�X���~�Χ�ޗ�WGS�JӖ��6x�\��{Tgk[�|�>|���Z:���=��Q��VF���o �8Zw�ߜ�5�p��d(��u�w ��}�X�����ƣ�w�29 �Y��P�������̫��	�5�yc�����j5=+�z�P
�w׵�j5
�ڮ�.T˗U���ա{���w��u ����!I�uN�/���vs�� �^Fj9���#2�?b���_��^���ho��S�V�"�,�����:��jHK�ZC:���5��N���Qt��M%��+IGI�=�偸��X�j�;Ϊ��?H��(�۲��`56��v���M`�ZenOz\��5�tY'�?g�>�?v�DB��<�j�yz<������F���`��$�Ȭ��Q������>s�j)�W`zB�������X�C4u�%��f���H�/�k����p�|��M �:��j)��we|*�V���� �&�R�g�5�T\S���)#ߖs^��w`���}1�Ϧ�5�K[����%ˌo\f�DL�;�|�ؐu�c�.����R�5�~������7-�6u�ǚ���ݥ���ͳ���bĸ�&!|Gs۲=a�1����g��'I�Ǩ��I�N��������vᆋ���v�#0����e�nN%u\��UGlj�T��R�B��iex�M%&޳KnE�P	�Z�2,n��Z%�	B�U��dZ�j3R�Y�����c���j)���/E*�k}{�j'ò�{w2�%憢9(��b w}uX����`dMu又D@�Co�?O� 4��|ZJ<پˉ{3�n7_,j9�Q�ȔᾊÊ�&�mg��K����IW��{��:��9�j5� (�۫u ��u����R]ր�j�X�r�!�Tj:�{}�Y��F�����5�O��})ThUSAYJ�L�(9k
���vX��3&��kJ�4�O:��]��kyn@*;��Xzȑs�G>c�~~�Aa�T-� r���{g�!Q�y��M�yQƵ���0]ݚ���Z�م}�)��]	�nD��zק�H��� 4FJ�R@���]�c�Oy�R"���י*IY��JH�ߞ���ycP�*H7FD}���RG��jw��WW�7=
��,u��lȦ�v�`����� �Iו\��S.\��s�.	�  w}uX����`dMu�D<��>�������a��r.� j��ݖmbX��ih�U�\y���RGz�X&��9̷����9�'e�v�y����}�x$Mw��yh�:R
#�}��u��e����.ğ��A���ާ�Ʈ���J�P�b<b_$�I\�T���܈.�Rcc4��]]��e�v����e���ոRG[偑5��ʬ��ʭ'�q�`
��Y����RGz߸��E=�,dC[;��yR�Fؤ��/�ъ*w�v�o�X�C�yfA��߅�+3+8�r<�����{F����j�8mbĕ+��N�O���k��k�b��{�W�þ�{Uv{Teo}y��1@u=��κ����������xY~�ee���'�ٺ��|�{2"�b��qyM�p}�n�3W�>�f�1�"�Dh��ה�[�\g'9R˥G�ٗ��dGUmn�"��*�c���$�K�X�ž�ɋ�y�;�l�%�P7ߖ�n9vdj.���Z�hu������|یf �5��k���ܥU"�E��ť4֦��&�9�|�$uΨ��Z�]^ ��`�w�̯#]:��b�ͼ_�_���[�j5׵k��k���/�E����w�HL.�F㸵�r��Z�u�X�$5���i��'��#�xl��rd�WY�w�`!q�=�C#PߞkGQ9���F���qj>�r^�̫��.�P��Zjk�P.�l��_�F͌Gz�����jG��Xœ���c���Yo���K����x�rx��z�Q�㶕4�.M�Vݞm-�n�q=<jk����a�v�ǷV9�s�[�5�q�g��^D���b[�ix��������۰`^��jtv������|O�����[�����s���}��Ϡ`�խ˓�B�S�i��5V�w���R�t<�af7�i/�����%;�4Щ�_}՘�5����Q�I��x| ��-���i��ĞbHxs�X�j�5�#���&GΠ�)��{��]O`�^�4\�IG����^(�\陦�1P��S����.���jFfK˻�y#js��5�hn	�݆@<R"���Ԑ���ƥ�˭%]ڛ��)./{�Q�{x�����SP}S�g��YSڲ�)�eB]�x�5��� ��w{�>]|F�Vf��\�1&�V5��"(���s�8��)sO�-g( ��G��+�K�O���Ob�ML��c,]ӝ��'kg�z�M�[)����Z�r  8BBN
)#�kX:��7�wnC�T��Z��9TeV���XdN���ZDC{�"���XNts����Y�Uf��
�|�ȹ5�V�M�V'C���hdze��,���dC���������$7�y���Ss�6o�e�v�tA������ڵ�]���uT�{I$�1=-	��No1>���wyy���7��{^���˕%�h��u�k�Z��={FG"󪳩�Ʒ�Z�$(�7���Qᗣ/-u�=�"�[�:l/rp�ODoz��vɱ��3\�c7y�y{u�t_gn�(��V�U�{���J�r98(�w{�@�{���H�7:��$��YF�n �-�ʷPJ�o��25[宣�v1��5@(����!Uz�j��*5ߵ`djz�U7���=s�kW~�Z�Z�$�w�BQe��r�u�g�n��Ē«��I��Bk�Lk��֢拾[��Wb�4Nz[�><<(�6��s=\TCP/Ϋ0j�������Ř�o6�|y}*Z�o��k$�%����73�g4C�fc^�;�/��.eog�����X����$}�/����4'�]G����H�Y=P�lk��"�lO��b���*�e�L]�{s��Ҙ?n�����A�@�V���u�nᙒ�Idw�w燺��pX��j:�W][�1=n��ĺ�>�>����R�q<:�6��:�ۜ�+�K��
�/Z�r��UiN�� �SqI�՞� J����CPz��˕sU34� �ۓ��P+}U� k|�2��x�2�{��9�U��qIߵjHk}w�xC�=���ۨ�g]�&\9T]V��H ���hd<��j�����wV��tr緗YfQ�zCpz�%����V�)7�[�$�}���+���1�F�h��tT�#��n/�d�}1c�9r�d�\Ӭ�8%�>��ݢ��������٭F7��3k��#�����to$՞�����YqIH g@53�YWr eS�v�������8�ӇoB����4W��H�����@N��#�;����]�LTH
�
��sr�T`dX��u���(\]����$+�">'��N'��Ǘ.b� g��b��R�%��.�`�ЫD�a���d�١K���p�NjXe߳�_�[�A�=z]`���̓�����)���Aب�^�VSϑ��X�����PtR�rbw$@%^N�D�(�T䲧����,*.�ꀍ11���c7v�3ڍy�G ���S�1�N�y�"��C�bQ�c�Y�QS�cE�\d�X�1@H;!��>>^�*�7����J,��9�,���S07�:�ol�Mn1f�h,�6�UQr.qS[0�c�b�d��Tͣv�G���*��5�᷺"wb��EN7nT�˅��|�-NH��|<�-����swT�Po�n��n4hg�u��0����0fy#"��
5���n�V�V�BYϊ�u��w4�t�����S��3��Q��aō��s]v��Zx�v;-ɹO�oqmXg��v5vԞ�srvN��+WN�ۙ�ل���*7���`7
E��1���l]m]sun���2ь�Q6�K��\\�c��{�n�6S��nwGP�(8cW��N�:˗�]�x��o˞��&���mn�Ra��u���u�ZO��y:��*nٞ��
I�:���1s֝���2����ض݋�:����ϝ�s��\+y�X��A��|w;�n~l�L�ݵ�[�vO��Q�rm�ooV+�[��Ɗm$Y�5�z�tgmqqr�q��[[Ö�������8e�r�x�M\<�
��]�����k��r�L�9���(�Թ�+����чRs�;p<�����2�e�\�i�f�J���2��T���p�v��s��Nuvxl������<n�� 퍳�Ч�]���wk�ُ5�ڭ��2�݃J�g�k�s�<��e;/X\g��7m[��Pö��`�]��juƻ;���:��i��f�)��^2��Ӎ�4at{]#է�<= 5t���UJ��Ilޱ���H�%�@�FJ�rE#2`���c[�����8gE��w>#��sś��h��<��YJe��@`�2,e|F�s#�N�p�',7!���b�A�f�7TJ��� X#6�4j=�F��|T^��Լ&��X֞�C~;��	�<x���8U79�o~�������|'b�&6�<A[>zP���!ma���4���ȩ��=p���0a:Pܢ��5�����T�5 ����ݣ���Ś5Ɣ�|%��/���w���x��xn��|޼W���HY�ε᪇�S��;[�5�XD����͵n )Awl�Ȃ"l �Y���mIf�-n�Iڏw!܌�}��-��_!�F,7q �K$��2�2�k��31`�-p�=�$ǝ��H��Ƒ4`��AJ��&Cyd;0�"�d�E�r]l�����|�ؠsl��I�Yo`˻n]ٍ�6�,s��7;�L�,����[�ވp�m����u�Z�3q�"����!����s*B�!'F6�][]�-�f]ɸ]s;��w��V�o7Z �M:�T�REG,�Ucʬ�m��KkRi k�y�7��Z�����w�R\�����,�ӹ���<X*��塐y�K�f��t�F ���*��R]֔�����j���� �u��[�u(���e塿�^r� �7�k��:�P��}�5N��a�Y��\�܈pb)[�I[婐}���'Aqw�"
KIJ�p���r��)Qn�$�kz�v&R�8���K���μ�5|�� L�o�[�Oz9Sd�T4�����?��t��kpsز6�OZ�l�[M���ō�6"�{Fo���R�K��}��?#�Da	 ׍%�:��Ȏ�}���R��{'���F�Kmg~����p�<Z�"�[�I[���3S��W2��%��"u߶�j	���b��w�:���I�M��*K|e��S4�):�I<X�塨>���mȧkO����n=v5ܹͩcGOd"�Ui��kF�V-kNЛ�M����Y&���{�$զj�u��C)W�@�����"����RC~���@(�xƯBMBj�����}ĜSK����ث�A���:�	X�r�u�/��EK�X�7�iU��{�zm�&��+1/��ˊ��.���$�{��<'o���u��jj��̤�Z�T�)î�.�.�I7�12���=��u�����P ��# �e"7��B-�볱�.��6Zfx�~.�t=t��a��Iǜk;�U�i)��,�V�Vx������꫅�uW���M�����b���5|��I������,�Ӹ��ʵ�3T����ɐ�2܀T}z3ڝܒ]Ԁ(�����I�/�� ��?�������T�
�w�K>��U�ېc�@�G�]-�v�g��8�v�n]t퍼՝�o��Ȁ>��� A�=J��$��-Q�r��E�jO^l�p
�W׵�j5��du�(�ח�폺������X�Kn�gIJ�w���6�V�K�4�S�C+IFַVF����uA��29 ��y�2�yxi�����`z�M��߾�GPz��W7V�<M�����*��<��	���F�貼�g'EZ�OC�H�ި���^��P�iѮ		.��Y�Kd��qm�*�ȳO+L7��T��fJѸ���n@!U�07�yX�P�����dr=��؟\��~K��?;�Ǜ���>=�1%pz7��)P['w�
�4�z��Mۀ�1{��[�	r�eMS,��"�::�4N:z�]��N��d���'Is�,յv�u�Na�Z�*�Hsx]���������Ľ���l:��"vx�m'gF���ė-��W��U�S1R�3d���e�!U�����I*���L[�䲫7K���m��<Qu����9���o9�%�3%L�;�Tk�Ձ��:�G ��>h���:�܀Tz�w�nᙓ2��P��'�Gpz�3
�Tb�%Mn8�4��k�=��Z9�����˳#P����"�w�{X�P��u�"j��UE^�VV�� z$����F���@�TG!��J_{���CB�[�S+� ����w�#�=r��@+��rQ�5����D�QJ�n�vX@�ctl��=�%�4�zԈ�IF�ߔ9��wfF��z�P�s�IV�Q�����)"e�/1��<��j�����f{rU�*�r�'��}E9�g%ΊL�
#���ւx���Z��n���# 2 '�
�*܀Tk�U��������R��w�4u��a������2��y7�fy�p������29 �s�U�L�wU�p|H�q���#Pwז��u�3SI�W��n�v�g��u
��n5����� u���Ϊ�Uku�])���=#;�KG%u��kr�-Yt�b�֜�ҁcZ���I���J�����	w��R����@¶]�ϻ/ؒ�,�[7ϵ�y����j�}`��8w��&Q�e^i��-¥��`	?"/c`|����Uk�bz��K��{:{���5��o`����u��׵U=��ù5^iT�%A�$u���j9 �{V�����w�]eU]h�P�ÿ=�7A��sF��-�'�DB�}{VF���U\�Wuwz����29Պ7�Un��U`djߖ:����;/�UN�w��@%���$�p�啎B��ą-Z��=]yK߲܀Tk~U���o��<b��pz��W�x]x�L�S+N�뺰�!��7ז:����3F��-�x�P��w��C3%�V��j�9�Q��FG'��uV�Q��VF���~T��̗ZG~	H��5��P��r'q��& ��ᢣ�҅$L�S�����:��-�?�F�Q�ɛQ�2��5����o}ަ�Q@����q��{��d�Ko+I|}�sM%�4�7�`j5�펣�={�a��о���/}����s�;0b�s��lg�{&ݤ�k:�Q���%斣p����=r�@���w ���G�N�ZyT]V��^���Ћ��~{���˄�U�^��S��(FSf�.�yZJw���y,k��V������:��_�(�zI�b��N@=�y(�C����MC�P)YϢ�ʹ�[��'���ʹ�y9�%�<F;��G�=󙆣P��r)^������9�j"n"��X�n���S:w�����q���S��q��/����l�+�Xe6�/d<Wv�@�8�����l�Ϭ{��~|w���j��Q]y�t=�8�3�����ŀ��5n�ܡ��}j�x˗��D���z�vզ��=�<�=�^oK��3[�"�Vs]߃��3�#�m`����PܨaaE:�s�4�j��~������B����ï����Ip�՟�j(5i�,����I7�6����D}��'�D.�w-Ȥ�jHs\�� ��:����&@<��Rkuk�J���hd��0�5 睓͓!.�;��1��ʰ25/��n:��Q�Ⱦ,F�����D��]eU]hơ�~��:��S�=��N��2�~�Y�����u��ț��䌰�b�u�X��q�>��O���qS�Jr�g�!e�����'������E�G�l@H�F� GP��$faʤ��IN���)��x~|���a~��)����G�ɚ����Cد��\��s��߾��M{�ߒ1�9���� ��oށ}7���,V��}��5&Vkq���ib��9��@�����~�ߒI�g9�-e�>v���߱.}�^_Y#E���h���*��B�*�������v4\����L��Dף�>�M�DRϱ��i%�O�}~X�O�y�N}m��/�<R=gP�)��C7�ʼ�w�~a�Fų����j�禝>ÕHl9����G�$bcM��s�ʇ�Q�F�\wpy{a�W&2��LC70�/�e�\�Gt�.�a6�q4�
܎
ru�^�ڗY˻f (_'�;=K@�P�ۜ��w�`�������~Iy�a��=�|Sx������`������+fx�߉λ5�=�����绶R�7���.�v��{M=����&X��S{�1���p�����]��Y���bQs�M�ё/ٲ�}�~�kY�o�it"��B�������8�Fd���9����h����G�� �Jhg3Ӻ	׼e����{�S��/5��,�M���T�z�����}'��b=����DI��с���W�����7�h�V�P��땶��nFP�u��!�{zL�Æ��@e�ՇڸƝ�A��\�v�� ��ڤ3+���`3\u�7M�Y���η��?��==�s����.�5�Sb���R�X�Cޚ��[��C��^���N/��b��}'4D\�4{�8@c�4�-J#.>�ԭhNh@�,��f���^��`)��1��:.�[_3`=�6v�ƍ�Y~��~�.���&���.�c����լ#V{�B�Y3�0���^�l^P�� � Kɉ|4A;�yu��Nd�-a���R�[+n�'D`E7pre|Ƃ��I$��Y
��&P��:�ՀTrp�F�Q���(�5^�_��@�)V��b��^{p�]!n��h?6�>�vc��Tk;�<u"�q��!�[�͗E���-��x��}��w�}�)赴o�=�ዽ/�y`* ���xK��W�]���D#�))��J=-�i\q'�ܴj�·����u5�aMC7�ܢ2C���ͩ��n��.���=z����So�7�����oDf[��,՜��g�խ��?,<�랙}w=Kk�q��R7�xi��.��Ԇ�ig�Y�Ul��~��8���m�Ǿf~֬�	.��Y�a�z�S�1�(	��}�U���go������������T�%��+,M<�Pj,�$�f����*a�m�?����Wx}#��c��M"Y�^�x|=��>(�
� �V�$ބ�u���������>?����z$�4}��	�W�?iM(���h��c���8vS�JD��oձ*n�]ַ�{5kr����;�dë��e_rV�.����>�;bf�A;B�DD
���!x}���6��!qmh�p�	O�Ac�3�n��Kt�1m���2�\2d@�!BI����[�Lp�X�kK'E����i15π%�D�&nw �*����S0R�XfQ�
��Z�۰���(H�πJ�3��}�W��C�1ɾ��}�lA�@�t����}[�b��n����d�	bU;���b�VЙ�1Z�r5�k�kk���M����@��y'i��qwOAӈI��US��n�Z.g�-��ymq&q�I�vC8;����K��W�۱��1��dqU��@^����7���v�Fͼ�5���%�����w\w������|	:�r�Y����N��C��j0��tD�����
��Evsh�iC�{��Ji3��}��X#��4$տ����>[�vMJ�ĤS�~����W�35p"4}��0�+>~Q�&"�+���=�0�Z�Y{33�����п�Z�*�UIF��Yq��u�n�$Y�/ �_Y�"�1
���T�"�`��D2ڪJ�C�2��p=���U�q�UO�O&x(�*��R�1�|-���r�L��gͱ�g��?��	�"�=2��~�����A��pG�&�,�-��L�؎_�L%V�#H�ЛN��@�UE��/�#>߽4eZ�LA��){TB��:�2�=3+��3�F���0`�4
L�U�u��H-��^���@&A�(������X�T����U|�(��d�m!CI���o��U<ޙ��
_h�L��BPKm�T�}3+uD%�
Bt�f���OsNvJ��7�z`�s��r]��kbt�Vc�wP.�7(���._�  ���(���2��`�Pp
j���dL�zb��T���z�Vw��BE*��TB��ڪY�L�\��-�Ǯ�'	J�-r0���"�Kaln�DeN�@,j�-���~>���6fW�x}�
�W
!��SPمQK=���U^H�T�b��w}�M7-�N�����Q�}/��2�ޙ���a�hUp�j��^�Lˇޡ��?U�V1��۾C2�I��B�o>��=+Nq����oM�}ٹo�#3KK�}5��QM(��RC��ex}�oUU��,6�#�}�n��~����c�3qӍ�X-p���鎒i�����߯��g�[�!)���2�:fU�����TWא#��k��.W�ӿU�4R|"mU%��x�~�{�3�!X�bxBi*�|����Ι�~�3?|�b�\��q�M�SK=���&U0�GT�J<iI��l��~�r��N&��t���U9��x
�n�9mj�<?'���bu$�C��6�w]�@�M���[N����=u�d7==��v0,Iu[r��BV�Q��l�e�^��6� t]qx/o���8�I/��ݮ-�ή"7oi�&=<lk��۫�3��+S����uj�� wF@�4Qf�&�U֐���(\���-��������"X��|��Q�� �y�LϻA2 �8�T���}]|�{=3+�G|��Ђ���RC��2�6g�ՙ"aS��Uz5���χ����3i��.��$Wg�HD�i�ߢ;�L3��̟_�e�g��2@i� C�dۋq<�6�}w�>a�ĸp�Sg93����'���&o�]""!D	>�������o{���A���F�������h�J#p�wn�Hu�����5֫�������vX�@EdD�>�TD�DM��+�夶�3
����EVDpS��]x{�Sm�js�}���cg��Dh����`��C�ӅUh#�}sYT}���؎ ,��[֟�� �q���j�*'&�-u�h�P �ң��W�^ﾙ��B��i�8 �Ug�3}����=�V/�L�6)��B�N���G3 �"�L�h��ͨ�}Q����83�vk���o���w*�I5T,�1��~r��=35c��a��W}g�:��Lʿ{��/$L�pOM"ER��J����^���!`���:)����p XugI�hkspv���E�nv!Û[�L�\�,p!���(��D�!DT��(�Q{Q��2�}=�«ݠ��JKmU����O��]�!xP�4�$�'L
߾��]J�陶}�ԯ)kW��.���q�X"Jw5|�)�G��q�\�{�n�i�����s�'7���H�� T��j�]T��*�K��*Y����)��BCo��߀��?�ߞU*ݠ/f�%�(�4e���n��"��N^xCw��Z=��>��u�胖5j�K�	��ſ}/"/�H,�)۷M�.����15� ]��3i�CH�E�	�^Z��8�%�;����M��N`��{��P|;=3~�D���c,�g`������@{OvH�4X��h�Vq�Nrp�B3�F}���o*��QFh�������PE^�w];�-g�4��Ku5+驉`�s��t�!��J�Iy&�}� �V� �����ޛt]2n� N��=�v�E�Y��8���	���S)8��G��ʘ�\�V���8��>�+�͡��׭1�EEȖ4˃Y:�"3��^z<M�M��hž.�������n���w�	�L��:�r��iJĕ��RP�T@��ᵒ��$&�i�]W���5����[��+�t��A��ƫ�_d�ÆD�\����A�a~���<�ں�;Ƶ�MP��|��[�f��Q7�B8�����H��X7���� ��÷�h���<�����ͥ/�튟�٠GuC���YGU��G���J17ٺ�=En�+�2�E�����=�gp�s���U�y��>F��>h��.j��y�����ɨ��K�#yu��K)T�����<n�N6@���M��ۏX�/�c��Fˈt-j����H�[�[�pn!�b��h��7Ge�X��r�-s����DWQ�'@��P�cxi2p�l�;nN�g�[/7����ɛ�9Җ,n�Ju�^-��Nӈ��:݌�ٞ�vL�V�M7+/V(�7\:����5kf�N�lFU�6�պy`���k�ݠ�,�m�Ѻ:���tL�R����W�7�j��;�������Ջ6.3ǹ�t�y�1ѽcv��b[��*�m��-�<�v��{GPr�]B!۷&��b�ZmA�%��+�ɮ-��p[pʚ^C��u\����m� �؜Ӟ��z;\�͈'e���w�h��ۯ@����{����l���Nv��AqYم1�Rx�G�kB]�g�΋�WR����u��6�q�ή{n�-϶)����;�cƉ��:'�m�\��ut���&.�;��<]ٗf܋o=������2�ۚ' ���Y��8x��Z^����k���a�"wV�;��d�!�2���^.�׵���$�2�=r;���۳v��jƕ�Nθ����:��\x�_lK`���g��L��:�M܄B;��R1"�"��ݨ��:�����EO���yɱ��/nx�is1Lg��zSӃ(�<RÆ��3���Z�cKۡ��g��*f�f>�?]�>�sD��q6�8�k � �nƣZxN@�ci��X&�\����Q���v����4�o
X"h�h���i��7�_C���SM��a�&�؃�kȆo��r�bI^]�S�=���,�S�q�+(��i�	�I�f�=��J�S����t�>��d{�`D��x�;C����K��F�7�N���t��7�t��fa�ۡ�MP��z={5��ȼ3�߂�� j5�9��>���3��PIg���w���5�5��4o�j�c��2�7�L�QøF��w��{Mq>��d���9cL�6�)K�L��த��F�ϝ�6�HmNY����Lݴ�+�5�{^Gۙ�f��&�thƛ���\�ƹ��� ��c� �u���V�w=容�^gwb��)T����̔Q�wW�!q�T�Rj��9Uݷ��n��vɣ��L�'+��T�R ��5���=pቬ��铺��6B
CJN�`q|$dI�R@d���3:���V>�!a��|��ٛΈ9���%6��؉⍦x6*c~dŦ{_�_L�*����SRMbgG߀fmV{��~IE�&����Z�(V��Q%����Ir���Q�j��2m���&� �. A��6�8)oBm8��*�Y�Y��
Ί��A3��/,`��yY�4neu�8�:6����F��.�4Y��"�+ �@��X���L�<πS���v!DL��ɊY���D_vL��0�����%|��xbk�0|�T/	�am)>���.{���2J�s3ؾn����u�h�Qu�f�5V�r���[mڵ��̭�������Dv��0Ҁ���a��C��w�L�_�~�U<���2\8H�T�j�He���V��u3�nz���0�"�B�sb����/��Htb�jm���}�O�a�f%��K�}��\O��M���ս��+3�e{TG}�o-L#c�k,�t�F��������9��F��g�������ug�vwN*���R� ��|��^qn��~ĵ7��3z#X/оI�*��;���͊2�����Q�}.��D�(�j��9�Y�<djXm@X|�O���X ~�UJ�Q	In�k�E:��������W��w���yA�n��Rf��@.n)�"sz�������̬�3�7=�2�5 ���e{:��� ���\�fW��*W��3�}�iR�!#C����ޮ��P]��e]���Us2����*�m]b|2�F�{������2��!)/ �F�Am�sK��3l7�1faw>�(���S]���{ʩ+-�=^s8�誧ݠ�/�EBb�c����Q�� �6��!?z_+�����AtL4nu	�*lFe;OoN�*n~�<��f5�A�t"���?g�˺y�9lG<�7�Rg�����\y�brq�=����6k9�*����wcc�m��\�ɲ�n�kjw�˃���V�0:-��9�ta��*n8l�p�uŧ'FǄ�q>-Ϯ�[�v3���y���2	"��m���2e�^A�FeY����\�M�++eQJ?���k��n���m\F�m^�{�	@l�(�}�+u3츎���X;}Ȉi@mUj���4��RO���ŲIl��g̀��Q����a����8��D7U�/B>���'ڙ��F|��xV9F8�T�DJ+pd�m�D������;7_������f	���-}��6�}�:��/u}�+�g&&�2�����V����t֜nxQDvm�6.$]��*��oÈ �'t�Q���_}k]������C�,'�I|ȓ~�L�-���o��32i ���!���{�2w:"�X Q��6�6S�0�nQ��G��r��o����/.>�?O� �M8�r��ڛ�D\pb��셭cz����~XE�\ϼ� �� �����!���}o��.�`��"�υ�:�$o��Y)�{�pO}[��O������6~��}��n�a��*{lBM�𱚶lLM�ʐ�F��o�u.V���ߚ��Q$�"TE �&c[�2�zm9�|��I�z3�l���Q_{�i�{����^_�O:�A�	�[k��U��E���� �R�����׾܁9�|O����y䡠�������^Ok�»��5 ���}��~�������`��6�@�<��#}�֫�V�������������:��جn>��Ai��7'z�OV*QV�*jK��Q(^�I��_f��j�A��<�py�CQ
Bv���]�+���EV/b�>]��&ܸ�pΆR�l�=�Nn����b��w��g6 �׀%�r g��4!�
`��< �a��g}���*�sm��
�>���F��z`�ۊ'ВdN|�ީ��ϛ����P}F�	xx����A��x_L������{�v���i�	�{���W��FU��}��<#7��n��v��ƣks��W&B�!0v�&�:5�s83z�m�Hq�ݭ�����8M��^<qLn�n��Sɪ2�;[Q�m��D�M��v���8�g�şksj�0��36��a6Nz�QF���2I�ѭjݮ����_�x��k%%��+&��x����<��b��e��\��p(�GS�RB�c��}�5�^��3���iZ��p5"����.���^�gϾX�)?E5G�b.�#G�*�t�1�$p��S�φ���\����GϮ�+��Nd�7�|)�}�����#��O���	%��$P�n	Unj���V�jyy��}���Du�<>����a5��>�zT:���,�����\��k,k`ȩ���.��,PZ��	��q�q7���;o�}�m�Mch֍�+F��~G<��^S��䡠���;���>�Y�	��_L�xBL
r�C9I�������s'<wܚ�	���x|3s*�W�Z�7}�^`�^D�Xۻ�N���ڽ�1�3��ե+�o��o9�^�~�^'w}���"!(�m�w��� �sg֙ꨰ �9�Yf0��r�߅�4����ɑ�ב�S6�Ǉ܄ >Y^��N6�j0�x�EWLY�����3#iՑ�m΢{�,ԗ�&��O7lƸ#�L�Ң��u=�����G�/cJ�8���i0#G`S�h�ڊ���3�o+pE��ݹ� '݇����{���Q�����Z�gMOo�172�JTT�ι�5�B�*��̧��ݨo^l�F�ܪٹ�}.���ow(;�0�z<����hhX���35E��at�"\l�H��Yr���ךfq�S�"��DA���l9N�c�e��'6-b�Iߢ#����hF4!���4v$aC��������t�΋��+��i#�g�k�w�Z�mi�3	�k�swa��L��C�5��ԭ�3Qz�Q�E4o:���e���d��⫍����0]0!6u'�M��G|�6gyR4!�Ż}x)b�e�s�v�Z�'.y�^Q��O��=���k��]�5�g+���>���XT�j"P��M/�	�0j�L��j��e�UdN����e�����7�wqy���Y5X�n��>u�5u�e}�˷Ż�6B .�Ith�VGN)�jظ<��_�(��m��(�sN��Y� �*�B��T���WEC!ٶ��sPD4�Uy�7��Я�/F�O���(���sѓ`����R�Z���Q�L hf�֦�0�)�?T]f��2�ii�P�E��Gf�ס�ůo5���ԓ�H�2�,ܔ�TA���=�U�cɏ��&CN*�{2��C�wT�u6횔���up-�"Y�Ea�ɉ3��#�5��Aq �|D�iI�ZIb��I�p��ww���0g� "H�H(H��L����ʚߞ6Sz��U���~�'3"={F�+�����a>��#i{w�5���F���&s�b�3����J��V�L*X K��G[v�S�)*��9Ͽ}k���C���k�l+�'�aܣ^~��Y������߾�B�im���UV��T���W��(^l��A��0�k(���ٌ͈7]{����4N�K���S��#a�Z����y:3y�63,�r�qld�y��E9���/r���1���I#"�#���f���W[���<�JW�����{TBUJ!_�[���Z��z�\3cZ�
+[��R�r�]p(��5̏��v ��|�*���*V���N���G�[�Q��F�4}�O^�K`���{}3+1��
w�^��w�i���h#�]�F�S���uT���M��n�+�Dx|�T�T[[[3+��5�M����F�z�0."��"�_Lm��Y��ewO=���y������ h �rB0�=�]lkp�Zzny�zH�n��v��۞���1�W=��[��S�ܾ.�y�d��E���z�S���S�z�۳���z����7`ۦ�b��X�0n�nc�� �&���uMO�������o,h�co�j�{_�.��]sף�3���b�g\�&��n�-�!ʜ4}�޹�j}���ņ�}m��z���J�+/@�w�2�t(�|7�l�D(Q��^��L�؎ 	~�0�|[UO5�.f���<��k��Ͼ~�MZ3P�l��5�/r�^�F'4~��֧>+��[����;[jW0U�Ŏ���U�p�<�f�̋���̫ײ�W���T����xR+���]���*Ǆ������;v�c{36s�f��7�iE��ɳk�ň���^_�����$XA�d!>��G��O�k�����ax�-?"�-ڥ�����4|�e�̭��&<���tk��`D+����ޗ�;��V���!5DQVY��ɓ\Üo>�z��t�E�"ƂJ�Ej�QdW����i2��� �=��kO���~�4Q�#-&���uF�����F�vp�y�a���){�BR\��v�3с���o��:�8���+rp_<y�d�pqev��.��=�6��/�H$IQI�Q��K�-ߦW����&q�d7W�"ř2{��Gﯜ�x�5,��H=�~���'ɵ����8}2�Z�´��\U�#��a,nR�F���쿏����. �-���6fG�ܡ|�ܜAp�*G������I^{�:�J|�	�'�-Wy3�}N���S�6��U�|�DU� ����f��DP��|*yOƁ���$D4O��Σrn\�����yX[�<�jTʈӋ�6��F�A�&4%,���'��ޅ*�aÂY�SJ��T���&U�֯z^��}�*�J3��U#��M�ec��/����t�'�����'�{�}3\�`�|�L���qW�'�n��� ���������DM[������Z-6&�{��1��:L/3����}�Ϻ�2}���^�(��|nT�~�5��K-���NS����obo�����k�s�<ኳ�6{�f��X6
R�p2�,%n��Y}n�pWMIoOn��c��
��V=[�]�q��ƥ��ɻ2���v3M�5�ɱ�-��k�O;�0����S"�'���p���x�N��m��ږy8�w��z|�I)41"RFcm<M7�ci���j� R�|��t�:n��e��p�뭨��NX煚����πj�o�c�@h�g��	�S��"M�M�m��z����=��'P�d�2�xc=�e�FI�]����D&Cp���̟ymvDo����)� �5�<��8�i7P�6"� �Ph�z �d�pp���]��`���9��� zq��\�m��q^k2���EmOvnk/���[�a��0�/��E�7���׵xC��BA�!$�R�1c�Ƃ@���3's�P�~^�ԯ.w�B�)�'|������T�y��ǉ�"8*�~�>z`�lA�d���tɟedB������� /b/�d�`~�"1	:X�$�I���B��A�S2��J�d��}U����GWL���Ͷ��N{��	TQ�z ��>j�wC�0��Č�\��������l�~��]pasc�4�*k�����1�N㛼�0�����m��W#����]q6�i�L���m��s�5�B��|�ޘ9�/���$`F� Z	���o~��fM�fwb��,� ���󞵵vւ��6�R���)-ll��6���k�}K����k0N��'� �6tJ�?�~��s_]
K��I���}/ڦ�Q��i�	��΀�}S�"Ky;�#��Ӹ3��;��33m�t>��{-}ST��u�3z.⧺)2j7~$��'野,%�������~����{����{������=3��F�g�0c[��z�T�p݁�OV?���l�R �\m��[�>�x�9i���_�&ZQU��{�%m�L��	�?Y��dB�O�	�B�${�y�{{T �4�u]���	|��z$́�vdM�L�P� �T�b�Z �ڪ^�D��ME����`W��D�ɻx2M�����	x(��`��r��*D�"����������s�����t��50���ȺO-Ғ��@�m��h�8S��FgyQ�
�����\�P�c%O^>�qPY�BV��m�:��f��ɃlM\8�
�9�Z]<�eӫB��'-
E6�$FlU�[7R�:q\�Tz�׺��g�s�C�L��/}c��q>��?��FmT�N��Υ�b`��j'L���Q�'ow#hF(6.j�R�!��8qG��)���ڟ�7��u2|(�>��-
�����=�!L�\�s��.��t���J�Wd4��Jo����Q�2�-E�y<�~2�J�����f�����
(NWp\Y��;���p����g��`���6�2�v��6����b:!X��̕�Y\"%�ޱ�~2CWg�H8��">�>]}�x�l��r�W��z�.(<vz�Qr`�������4x�c�[
am(��.�g��bN�
�H��z�*r��<��9��az�x۵쯎�$6���k/I���q�x�_]�O�g�s��/ńݑ�wl������<�t]m�ݩc\ܙ՜�r�w^�p�K��u/�Ñ���6�Ɛ_^�˞�Юuz�����0�-֝�>���96NKeN�b綯�]t�����]rp;\\m��&���s=S��k�6*#mt۱�ɪB�p�e�Ų�ц��^5��˶շ*nNƬV�z�s�3��r9���q��9+���d�����Ǵ⸍���;�M�Mɢ����Zm�:��<�<��=�*pZ�vL��]�k�{�]s�m3��0������\��C�GUv��9�bkؐ�y�i.$J燠@z#8Ã`��s��SǴ��le۳;	����1�Wd7N��[���e�2��.��[Dpc�����&�'o	rU��k���sݹ�=��Z5��iw=t�)ȏ[&y���Р19*�EjT��*�BA,B����2G��V\&��3l�8�L��v�8gz��źz��O<�CS���5��pDlQ��;j�ۖw��9h�mnT����y��~��{v����h���`��X��t,��%In��C	`T�/��o^9�Z�R�Oj��(f���s4�L�E��%�0iY��^v�
�Dp�I� r���=�Ӆ��Yڍ��b4;6஡@�u�oM��lOqo`9�ë	�^�#�`�C&`p>��s|��W����3�������6w.�>�7|�� _r˚6��cP�ա�"�|ǡX�������K1l-U�9u��I�5�]�q/i{�{+G
�_n<@�{�w� �=~ �b�)
���j���"��Y�K���˞����3EXg�Ktwg��v��z��R�
���ϧ�%�>+"�K]F^Wt�]N�u�
��:Yȸ��ꗷ���'A�4��n�-�3���s���u����[��-��� R�*��r�Ѽu���k\q�i�u�ջ�y�c����7�ۯ\ta�ka�(��Epݻl�`5Zι�vgu����5b�N�StW[�J�_�`��$dDM��뼞�����bm�������<��k��R���۞��֞�m�������s����{�օl�o[�����癆_Hmcmw��|2�=��mKj:��)���p]�e{=f�d�A�Ȫ�O�5Y�&W�>�����8��Y�*���^ ntѭa�M��\AR��Î�w	�1����s��{j�*�ڋU�.�P��&��[g{-�G~��C�ٙZ9�L/D�N�ksУ��yU�м
%�jT�����)'�W>��hm嚾;�НZq�:���<������4H3CD�)b��D+W��g��}�͋�My�&��+jj�pO��Fu��Q?T���� #�޷+z"%�Ώ�f�4~�Bބ�U4�=g� d�7Wt�Z>��	���躌� �bƸzQ�Z]$�̪�5G9�t��I�[�&^�D��i=P���8J�#�):�i���"_�N��?�<T�~e(5Kz"VD�-q~�u�&a�c�ķbkj[���!��S]V늫o�tl�N�����=�R�`�bm������m���M�<��i��_~K��?l�ج��:߇���!n����c�Y3��B�X"��Dؖ�q�S����}m��}���mBOd��K-c��V��T���d
6fɊf6����|�U����|)V0�^�gC����ޟ�I{���!).���p��ۂ\+"i��$Ͱ� �far�(�����HTW �~�r����D^�iQC "f��;j�j�F?38ZY�q�*ڛ� �+p&q�}�EMd���G�23> �H ��$��!0�H��55��k̼ɕpU+xb���r��^��|�x���}3r����=�4�;*���B�Z����m��n��/,V�l&������dD7����j���8�kי�Z6��VAO�ba�Z�iIx PO{��舡V%��WȔ�V�guL/�"!Oz$Ώ��
��#D2�5H��1+�෥̺�����Q
��U�.}dVl�*;uk��j�����GSE�W.{���}��%�v;m�MD#ƍ�P��K���:�x�9.;mtT�8��sqb76|�;K�z�ɛ�2k�r���OgO�v9�]��'�f��r�=���t�s�������s�ӄY����Q�����uc�uEt?~8�w��5�b�r]{z��g��[�;7ev�t��:���\���aT��ks�޺z��*=��B(�tĭCy�|ʩ�}�|>��Q
�"�D��^���#ÁT�ѻ����ޘ�}�eu�){2�:������,��3l7�a�Da���{�I�Z7ssﭿ�N_z]���7�l�g�<u�7���#�f�	v��7i�v�H����-pq��	6�?~�_l�'��V�x�EÅ*�~�w�/6�(��ԙ�w{�2����:h^,���D��N���$M������q�|=*�_j�&2�؋
`����׮��ؓ6���C}��x�Q٪Z���c|�t�rٿ�����K^ŭ��^��|z��SN�f`�{��G�~�).��ݖ���)�~��=�'��F�d�C͕�ځ7n^��.XF�'��i�A�ȻX��+Y��{���2��B��n�QªY��f��5fr�$�0�M;�����8�}lA!���y5��#��������t��2$�&m���@K����L�w{�%V��O���>��_�et��b��o��}�l����l������Vɶ˽.p|���--��j�_�!h�2��f�m`����"
�dY���x�:�krz��ϻ^P�4�6E���R���K�	�^��~�af��U4��~�HrJk5���R�3�'����(����u�U�g�sI�e*��,���{t�=���ܺ^�T'Ka��VD3
���n��:�(��ro���b�j*u���}F�wL���ZJɤ�ɩ������/`�T:����f�c�E�`��#�߳�3�Gيx mٹ����m��6��*��������Kg������?}���(Cos��,�����I���	��J���Q
UK=|�ٚ�}ϮާXI�q(Yl�{�a��ѕ���)����\9�}њ� ����$������wD�^N������H�v�����zԋ��%P�q[9z�7딣���0����C%��@�`˓�B�A8w3n�mS��t��9^�&�%�7';kGg���Q�EF��Ńn8�؅�tvTɣ����8H:q���cn�ⴞ:����J�R3;:�k]{l.��5��x=�$VI E0ªcuV�����l'6�՛�4j�%�e�4"c˵D)�럀��]�>���qfMk����rN��԰|8K��n�Q�V��s�:��m�>(o�m"ܬ-�3���7`}ﯦM�Q����n��GG���R�#�o@���`/���N��nz��n3r<A1���4�@A5g<�
�����������
�9z!���L=97����^67�S��}wD�=[y*���s��S��[��le�39
y}����ȁ"�� ���kus]_kރM��i\�o�d�\ Qp�k�R�^`�Awv>��Ro[�7�@�>��NC��Mk| �y(����Q~=�=���=q]as:���llQQj� Zƣ�߾�w��"�J�Np�� �9G���^�W苗}3�e����"��{��M��y���<��9U��%}j|6v\�M��c]�-,hbD�������s��1Ln���˞U՘�����.c&v�	) �����`<|����� ����mm�c��mFMH�C{ki6Z��ܽ��p�V�[��7���T^�%��)LI���j�l+���x%��5m'$���A���O	3�d �:-�6x!��v����J.�=��S8����o�[����]J�����`�����EcۓH��,��˜�?.�'����	Q�zSv,[�����2{��]��*��p���2��i+����8G�"�S�Oi��#�l]�E�����y�=�o����g�����{cU���)�<�)�M8��qښ��;9�4����&�\",����S�v��-��(V�)7�Qg��5X�ޙ����Kf��yT@Hu7�e��{���fj ��
�p��X�S�/o��gyZz���0��v'|�wN�w%ݚ�p��"E(1# ��AX$o�W�C��DIM�?Q��3s�)�R��e�?_bd�7g�6q��tr���� b5�43V-x ��cX������8�|��{�d��wA�vQ�4@�wEi�����N4�/E��+96N��G'�t��ӦW�u�>+Ӂ�vdəq�v�N+�B�N�k�#l0U�cH��Q���}@�sN�˓����(MU�Έ�-�/�����1���Vi��)���1�\�U��NxQ���3�^����,�4�!EsB���-@��հ�'��H�0L����M9��rS�e[�(�n�ҩ�����oN�p��y@�� ��o������,ش�;�Z�9�w !K�熫�5�K8��f'޾i�E5U��'yM��_W�ua�P���s8�+@��(MO��,�}y��;�� (KsC��D$j���� }�3�ڠכ�>&�,BJ>h/��s���:)��,�_�o��b
'���u��7WB7��6�p��^�ﬀ6�5������: ^���n&ER\[Un��{���PhP<|��)߇�7�2���=K���;��n�
R�]�Kj��$��:�:��11��N��s���7�i�E`I#�֣Z�lje�-�����w˾ND! �@�ky�CDem�7͙��Ջظ�:��GZh��B�[�XuF�Ux�\�g�����2Q�{����}`�P���ԛ�
�":���}�Q"���
s��Y�;(N�'h-��p�:$��*�
������#m��+&���v̼&^̳�s[Gv��ې�r"Ue���徻��dE�u"�m!0:�jΎGwخl�B��5�:�E��`�����-�0�LT�ڝ�lwcq=�]ה1Om�s��m�.��-ɮ�s[�����7k�<��Wnv����m�<sLַ�ƺnڷ7<�]v�xn^�Tt�n�ٕwyoJ��D�ȃ"����Ay~z}�j�U.wbI�R�l�����=lG���i3�Ȩ�K�aɾ��霽pqL��|�`/�Cl&�3�ٹO>��t3[���f0�!9���󥇍N�Mb�"�0R�~M\uoE��|$Gƴ�p�q�n��n�ƌ���z�n�`WFZRM��z�^���=���2�z�ҕ�s{ME�u��v�sx��yS�kN�c*�\�
Ea��׻)p��S�n��O\���o�U�[c>YGR�'uP�ʓ]xxu�^�ՇA�;��f�}
��:�B��p!g@�_�K'->���ډT/O�"��T�ޙ����^�k�j���Ln�o籎���:����X�t�q�NQ�냶�HIÓ�����U���*���eh���y�M�R��>��Ř����� ���*G�UK}
�&}y`���-m�g�Wۊa;�Cl�<_m�IK�ɾ3?*�.*pЅ{�������g�� ��E�[�{��ٹ�{|zU���f#ﵫ;�au(� ;�Dx�G8�u4��ҧ�|y�4q���YԒ����G<B��9Z�gHt�Yi��I`�w6�TB���^��T��ҧ�ursm::W�ko����h}��>�{r�f{~EN�_#�:����^��}��D=3l�9����)�+�g����ەƸm�gsM��j݉�z<ڞ����F8mck{6:�b4Р �H���qG�Rmz��{��IKl{<�Y���Ƿ8�6��[�8�"�XGqG"�+�Tv����EhE-��-u���_%���y�|������g��h�]���6��ݖ�Pʎ��w�b)��Ե��7s履j�x�������3Vt�Bg�x�-u�;*���8�b������nI�Ю�cMok��B���_}��
���jsp!��)qj��9���p���6v�]�N1�a�6�h��=��v��u�f���V���չ�!�G1vlx�sļ��8y��{x���v�Qۛ�>�P��ĝy�������.���U�坹7������,# 5G&�Ce�1����L�%��.��Kq�
`�l]r�E8f&��dY jd++D!4��=�������h ���W��Nx���7�mzA����%5|��j�#���K�12h��a�T����ȏ/Z�^o>��12���F+�S�^�2�T�����fAnCp��w�q#\�͛�C��y{TȟFv�����wV.��~�s3��	�iI���}q3�Df������^��ߊ�*yß< f�$��������O7�5�w���۪�$A��9�/߾��&c�{_"�|=��O�s�L��9Vfi~�K��t�{b#�	�*ߌBU��V���0Gǿ6=����=6��q�b�0����p�_G��˧�b�Ep���s͸̲=d�a���?߀R]湕��I�`= C}y�C��g}.dD��,���H�ɬ��ӯN��q6�u5������ї��<�W]�9�$�N�T	O*�9Y�[>?;g�v��쁭��L��]�xA)F"�k:\#~�̶a�5�B�#�5IW��W��&{��/�?�@!��Yp�c�]�.Y�Ѳ�. �혆ȻX��#����$���2�dވE8d��K7��@��:$ΰڇF,2 ����>f$NE_����c����J�ʠ,za�C	��tk��.��K���/�D��wR&�u�r���� ��y�3�������L��9�&���νŉ��fԜ�'b#(N2Q)����B��5�/g�L��f����p���:�*��n��̷�se�(c����»��?Z�����~1�#��n���]|�&o���l}�{�]���L���?r�X��|��y�2���3�8��D���<\f͇��߷��WkoO�O_��%��2�۝4k[j��P>=2�0/�%�E.��g�b��
ǘS��>+��H/u?)��{���@���P�=_I�ɼx���]�(�0�A/_��S�QC���y���dWr�#�;N���W�Y�����?���Od{j�zF���6�9�v�va7�7ګ������%ϯP��*U�Uk&W3�vj�*�n�&֊͈{��s<�G�|�^��])o;&(<|3�sS��Ѩ~]�1�?-����G���d��5�������=�g�~��"�c]]4;;����L����mu���^����v"�cw��ym<�j$��R�������?�z�r��<��
gM[�oT�^�y�#�e^�a����t�\�:/��|]\��ud�sh�Hc��^����Z�<}�:OEg�tUd�;�֡C��u��]�Fi�p���)EW��������c�:�f{aR�~�㴘&py3K|>;d��2��s�  ��c+lD(�ڀt�q�uتfݎ}��lm�y���=�[g�ؼ���e�FY㹞LS-y�.-����Z?s|���{1yr��d���]�$�շ4�<����i5�C����lv��j�j�IIm]m���Έ��q�7N;�g�nB�<qȘ��vyq=��$���;b���v�\�g	��N��kX����Qd8^�����/�s��۠��
�����vڮ��;�����7q�
6�i��ܖ��Z��#7ma�r��v����[�{g�p9���y�&�;>����nZ7�]�3k��=�k���C�랢Z�*펣���l0'��]�hω�Y�s�<��2o);��;rb���C�K���\I��:��sS�����h�]س]g�n-���9wFv6�ۑ��i}cv鷪M�����97n��=ec���;�m�~��L�oU�e�A݁3(�A۲e�8x���8�vI�vK�8�� �v���2���q��5e�n��i�]#�2r���4[{Ep����Y��Ӯ$�ۛ��=���u���-;6��m��y��8��䳭�=�(�k���[�9��g���A���?������H�Ռe�E�9[Y��e�\U[�m�k�F>�Z�� (�|��z}��0Ff]xy,E�ZJ�/�� ���U���SL`�iR�)�O"�C�(_�ደ&1 i9D��Y1�� Vj��	$�!d2)]j�]"�v��<�ެBo�6'��]�J�7V����WS器I�i�?A�7z��������HÜ8R�d&(7 �~��XBt���v�,�i2`�ɑ�h�a�B������y���"��:t@�J+2o[�։4�]�Z�M6����W%�y1�8֘��x554�0��(f<y5��z�&D��8�KI��M����Y��< �CI�N,^��3���N$RF�3Ma���ċq}FR/$�F���4�;����i��BMu=)���$��;no:�w���q����׋gU�]m�����\�,����yݬ��H�2�{pp'�)�����mv{P��y1��%�㪷#נn��ǌ7:g��Z��g\�75k�9�[���w wx���7��m'�۪M�b�E!Zd��Z8{\񧌒�Y4|��/�A��������{�ec�� }2��9�s��4b"!E��|c�.�@�6z�4}����Y 0�UK�������>���ԧ[iu]�b6j���[�p�6fWZ���O������j(�4��ҽD|6-�8폿�gR_~�k�V��aO]�˲:�nM�^/����☆ଌ^��шK��~|I~��Sx#�&ϛ5�+zc�z�\+�ks�)Ԓ8}z���6&��e��E���Oy;�خ�$��y1T��s*�hw�U����>2$Y$I���ߺ֫��8$u}w&}��Q���>�[9���K��4q�4�c��T�@��S+�D+� o�L+c^q�H�J��k��b��>�p��ft��
� ���m�$KG�����K�]f��;����5v�`D%x����������3!�d�j�����y�3+�D+��|%����[�
ib�Q�7��rذip�Q�5�s��Fs�=�&�f�s���K���h��I���I ��?��}�C�T��`�n����*��BW�������'#D" U+~1��f�_��3��S���1�4��������֑�`�ѐ�Z�(딭²cr�rO�Kf�l���/�B��ܒ��[�K����Ulw)��BW�~�e�<� ��U��Ɍ3 	g�.gL��!�H���5U�|�4��y�!W�����ߺ3��N��9��3yK��KatV ��&�#+��LN�i�s�2 � ��ȁ���6�6�I�7�	F�k�����|36g�ڠ߮#x�1|p�'~0�0T$��)�ɧ5=gd:��Lj(�'پ�ċ��Bdv�n}��)�n
�>�?}��{sɟO�w��0�~h���X��(����>�85gW�	����]�+rg�h�)���p�f$ʖ}����y��97{�1�e��"#�e�39�=X�����W���	�'���.g{��1Ƀ�9@���H.Q0�u�Wjǝ��Ϯ�����𛝍�)&����;������j�5<��Gh������m�.O�G�飂�07$�e��Y���ݙkv�򮩹�T��XKK��g{�����c�M���%nځ$�m0�V����:�m�b��ݹ�&�$�s�H�T@�>�������2W�A5'=��%�}~��|�}�P(]��A�Iu^<ѻ��>�ؙ����A�|r�N�'���s�#Qџ=�n���jg����>�g���>���v#���O]��p��Y�m�����+u� N�<�U��?{�x�G�_���L�ؠ��+����G�Z#����=�=�QS�9vÌ�rx��
�򚽞s�:����w�~�u�FE@�d�*"" �)eg��{ߔT��t&��眢�a��w�en'<W0{�<.�Ђ,DD(�߾a����� �:b���DB��Rs����P}^ɟ ����-~��U��t�vGkv�Ʈ*����J��]�9��M)�wU�����/�xa]�$�'��|k��Gx>����>a&!8*��/���q���ˋQ��?��C�����@���NEWQ�r;.�`�CQ������A�]"�ڍ�W6Ŵm㘕t�w�f��a������kaB��ftڠ�YЌ8D�Q������*��1�l̬�<H�C-��p~,��)��ȖG4�St�H�脃V�ozfy������Bd�F��!k�|�)�_0���������}>�pIK� ���؃�hz}u<�,H�-���!X>�Q�؃�c��Y�~��z^;^܀�� @���Y��djԞi���$�e>��z�3�D�)\��0����+kh5��5\���Z-�ܷ4Tb���O]��#����t����>���=OusY�.��?9]n����-*!$N��*:8:Ie���ܡ���מ�rpY���y�xd����}��P��FO���Em��`�Q#�3��i�B���%������YO H�U^�pb!1;�����'���Dlǯ�f�~�&vQÞ�p�Q�j�Y�ǀV��R��w�퓽[ʐ��wB,��}�����4���bEջe��=��u�^Ny&��0�8㫳�8�'s%�I�j���%a�ɧ���r��Un��-�u�m:ӂ�nE9u����q���@�{��ݻ\�_;���73��>�4�`�qlh"b*�oq(�X�۵kE�-E��b��o+�ޱ�CyKb����p��q��e�6�p�N�k�k}�b�_����yE^�j�篟}��6"�b-Qy�
�ݿB����E���ު���Wo�I�N
�gt^[�x�x��揳4��.�+ѵ} e���-�!��uv�uv����bp�j" P���jw�
 �Uؼ>~-A��U|r)���d�t�25��R��dV�9�7{&�1�T)�q#��GK�.�ڛ��x�)�^B@�H�m���Q[sm�f��*ȡ"�� ����o�	w��Q��$bw���ь�x���<�H6,���N�@z`�(�z_�oDb��D2�s��w�^��}��}��`g�C�n�vq$�PN�����hb	��.v͜��E�~�G��+��	�o�%%�n}�}^xY>(�z,|�7��&""�����ؘ�=�1������1TLe�fH�K�����" 0���Hy4Ǒ���]��2l�1(\�Ѭ��Ǜ������1�.���DA��H�}͚	�����{�^�H=�+��U'E�h֕OM�ϋ�T�ǰ�ta�A4)�ɐa�V����w�.:*�`��.�9��"�LȠ�v�5z�f�M��������ݥY��AG�kUf�P�:_1l鿅�ߌ3�Ud�ظJk���C\�.���Nr���=7ӚNq{I�X��V��&�~A�Zs7w:���_{Bw�ޣ��pS���u�n��L�.Z얅+�T_d�w��C�?,�#E���ojej���o�N6�+�D�3৷yq�~��c즸�B�1����裰1Ă�NVźmMȍ�h�1C1q��,Z4�ec"6�/.ܢE[�D�#$]�a��:����S���N��R�g*��HsH7�{�u���O]����o���<J��w*��wnOQ�s���/T($�T�x�Ŝ(�Dގ��zG�T�֬յ.w�%9-�
�גaEb���RI��-�}BL5LZ���X�5ơ2���U��-'�ޠ�rk.>�U�m:$7�#)����M��#9F�c�g�<s;NT�r��ڐ0��Xvh��r��(U�Cl|�ˉa9�%1�������1�1�j��Nkۄf�!a��}`_%j�\KG	�N��1�D�E���ek����p�j��k���T�w����e>B����peѹp�hӏ��E�j^6��m�j�r)Q��<��8b�88���5��`aM�����3�bcm6�mB�dͦ�Ijn�#V��i!��"f�l�R��X��3Ơ��	����Ԟ<[�:hI&ɴ���'²e� �["�lc]�Q4��a�qͿZn���Ƥ��M�ey,�b!����UE��5xڊֹU�U#�
#q@	�������S��\r�=U�ex���uʯ��%{v�hw���6�Q�7�{�Gؙ<u�>��/�����٢��dVx֨��ج��[b���{����~�	�G��c��"\(pӪ>��������H��_	P�[(������7�z��'ؙ��ϡD*&� �ޑ����Q>�!�����aK�����޳��L�QT���L��x�| ��wkx�ܶ-�F�ض��U�E��b����&�W����D����fOgtπ�A9���s���m�q�2G]RH�uq�3tkzy�,Y�//3���ό��7�}����fo<a7��-I;��)����&,�Ǒ��HB�=��&t�'>��)��/(� ������`��#~�,�~�pbK��S��6{�j���#��7_[zI]�3�va��ёΓ��Z���u���̣�0�oq���+��S�C�(��`�H�F:��c��F�S���onޭ��N=��z懩m�{.q�xͱ��u�ƒ��	]@��a8�O嵰5@j9xN3�:��dg����89���NvѦ��<��ɉ�3�){]OIsƛo^�z�}��kc���V6��nV*-�j�͹�����5�N�qi)�]n)kN1��%��J�g���E�t�3�'��yo����W��l������F���d �R�:0{��R��)'�tϭ��k<���>�EXLDUh=d�tA�7�_���RQ�!�&�����w�Z�=4���{?7��Ev�+�R�dqvg:���o�n��m�m?a�7u�3�|>�,� �b�B�1j���O��l��7�������;X�ÐjN���-���9�7��\�����A{�TBA��U㮱�[�+��W�5<m��ԑa��_��~�0�_��#e��>���#�C�,mq��\������x�z�>��*�s�Q�W������?~�Ԓ���ޅ�j j%jR%hQ^0b�5Hݧ�g�x����e!����=��O��l?57�~ ��S���
�0���-w�Z������یU�hW�"����7����ļgy�sn�jځW}y��؝�p�F}�XT�W�}5x�n�ݷwsp+s�sb�m�oMs�tt�Ҽ!�����"&!O���;���Y���·�B��|�LX����tA�؈�غ���S��j�J�\M�*('S�ܵG+n��r'I*"�ϽBo>���HS��Vz4ZfN{�0ҳ[�Ȏ�� �x�8q�^��߇��'{b	d�����ﯶg��}��=��.O� G}� ����'�x�3wuM&��{.+(�v	�ˬ2��^є$�󺾵5�v�# Ȅ�'*��N��gs�뻑u����o�=�g�"">��z`��m�!K<�u�o�hN>���K۠��K�x�9�u���E���Z�ZK�������8L�v`Փ��ЋuG}� L��G��+�o�J�=	Ke	�7��|����s'���.4UV��u;��!c���-�l'!C#ڷ�V�{#������fb���61b=�gb�T�i2��O'�˹ x����'��S.��?�����9�P�+ֹ.���\�#�\t�v�y1�8XkЫ͑�i&c.�{dro,�槗��m�3��Ⰹg���:{nX�g�����v	�NK.����h���s6-]V�)f�����ut�E;��'�{��^�'vnG4�+��y��|z�^;���\u�8�.��x���;����]+ܛ>葾��m�Y���[9Ç�6\
�w�=� �p��&}�3�0�~h�g�7�����w�f��`�E��]�����}G﫦��{����z}���w�l��g�p�l}����<.M �X�E��@�%MZK����\v`���+��xX�|�d�U�o���{-��<��Ts���F�:�����έn��b�0Dޒ,�TV����\�P'gw��o��oȨ�G�[�r�!���9�A�q���fY��(���̟sfj�>O��S�١d�7���U� ��^kq�F,�l2D�>%c!����?%����?���f{���蜉�yVL�b�3-n��M�f�<7t}""����N�fk� ;��q�?%
$�y{��,X_y���2g�v��%	����Ϸ��@�Ļ�+k�lFgmB��b>����q��DtL�C�*�7�ۯ�z~���%>���bQ���NLoM�����m��e%l$z��wDN;0o��T{�̄�Æ�� �T�/^o �[����O�hq��ɴvJG�i�:���@�U�&�>�k�;o>��fo~�<��	�tڣ�? b��^�{ct�Ou��p`(*'����o�*w��a���0�0٪߀��Rk: ��#�>�D{�G]���/~�[���&��U�N)��b"К���F���%�U��`�ڦ������}��=��Q@*!r@f�NM��6�~�Rmg(>6_��ԦU���{�Ϸ�ݷm�A�YN��)F<]���eK���1�����1��3��}
��C� Bj0��}��yj{�_h��<5��[`�U�S}�K5>�G>7b����l&������_��=�܈9��9��Q
��þ=E�k[�K��?��'���#'� M�[mS�~�km�W�?j��@���?�.e��QE
�kM?��3F �QV�*��V�m���Ű�5�+k�����64V-���b�0U�UȂ��Q�P kX���T[X� ѴF�
-A����d��(�DcDA`*��b�E��V#X���1mE�lX�Ŷ�b�k��ETh�X��m��V6�4m�m��jƵ�j5��6�բ��U��n[k�V+U��k����mlmh6���nj�Q�b�5�6#h-m�EU�Z�I[r�Z�*�h�Z6�Tj�����[hբ�ՋElU�Z��F�j�[j��V�M�����D�a TB��ɬV�ѴZ�M[�-cQj���ڣ�EQZ�-[��EF(�WM�{|q�ѭ��ccE�X�ZصEF��Z�FѶ*����"�
,F��DA�"��`�Z�ʮX�j+lch�kF�*���Z�5�j���ŭQV�kk���[VMVMkI��%���ڲ���IksXѱ�m�V�¼���kXڱ�1�����ࠠ�-Q�b�b��\�X�j�W ��"�b�
�[h�lZ�mtڷ6�6�(**�F�V*���V+h�[@[h�VD�"��lZ"�T��P�d@M�!� �FɲUI��I�)ZKl�ou�򴖒��i-Ya EQ�/t*%��\�QdT�&*�� �"�QE�(�dE".DJ a ;�dN��-����!�y��'̥ dEAa�?]5�u�nO�.��ӽ�}�ϭ�o���iO���_��_���t İ���>�����?��o�z;X[��?��X����}>�t��?���DP?$�b�����i�?�!������*��?Je�@��c���>�����~�iO��>
(|�����{���~G�DP �"����v/��� ���h?��LH%�k�m��F��ޱ��Rֵ�����������O����
%��g����~�RE�A$Q ��kF��6����ͭ)k3k5)�Jkif֚��"�H�@b�"��D@��H�A�$A�D��`) `�")"�")"� b��@V(��$E`�B(�"�(���mimJ���l���kjR�JV��U�V����EB
T �H��B(P����@�1�)(���5f�*�)�(�EF�J�ыQE��M%�(�k6�QQF��ղ��Y��ԕJjMMkfc�U33i�֘�5���Ym�Q�2ڲ�kJ՛lVZ����-ka�Ѭjml�Tj�5��RjJ-�VTEJ5l�e2��S[MQk6�I%�đ��([Z��kk-�jԪ
��B  �
"A +H��A"��R*$Q"DR*Q ) H�E 1�Q"�H
D�)H��D�$Q"�"!H DR�D����Z������֛5�*�kM5e�kE����6�U�-�[&֓kL�ѭ���6�e�ki6��m,��Z��Қ�YkJm6���6����S[J�ZZmi����[5e���Ք�ږ�֚�kJ���jmiVmi�kiT���kJ�ZY���ZSkMMm)��5��U,����em56��Zjmi��"�,Q"�)H$Q��ʔ������YMe5��)�Sl��������)�if��%%���aR�"F(��$��MZT�ҩ����6�5����f���6�ٵ�E ��~(dR�Zy]0z [��&������P�(�b"�A"����}����8�C� ��w��*�<�>��4'�(x0s���c�8���寡DP-�Ф��0~G�~����0���B&ڗ�s}��'�X�??<?w�~��~z`P�������>��u�?����"�~�U��O��X�������?d=�GK��}�󀊀�忙@���?�X'�4�kq~����E�~A���=��p`|�AP4i�Å!ÙEP<
��!�S@hw���J��Z�����:J	�p�"����!�O���'�g�@�F��ȿ��C� '�.�����|}��>e$~K���C�������~�����O�(�����cݪ���,b�{��̈
�|�Ҋn��~N>�����������"G��(IKl��z'��c�/��/�$���5��!����T=��� *���PsYT�MS��G�" ,���@XtN����{E� �M���c�?��M"}_Ї�>�(���4?�?5�E?�z�ߗ�D��*��'�P�������t�Q����^���Ώ���3�W����.�p�!'@�