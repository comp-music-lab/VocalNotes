BZh91AY&SY��l|�;_�pp����� ����b(� 4     (                               �            @                         {��@  )I
E@%@P�T ($�UH� J�
 �P@��B�BU$� �       �  @8 |�\�f�}����7ˮ����}������=��k�����o6�f獩����m���e��Nn��׶�ۨ�R
��)U"� P}�WŪa�b�����)J���]��J_-E���K�R�������t�*��{��T�k���yeO����唪SϪ%	
�A^       �����7ԥ)e���ꔼ�����W�R���q��U)y������R�Y|o�#�)xxwJ^Z��Ǉt�e� xFU�_Ox�|���
6�HD � ���J�Z��7OJ�<n #ΕB�^}|{�)�4xx�)��U{�|�_-J^���;ҪS3^7�UK�G�����*>�󏝟B_BR�P��      �� @p �="M�t�^m+��/3J��&�Jxp y�J{��ҕyjW��y�uU�}�|ޥJ�. ;�˩J���=�<C^�J U�
 �ک�ԥ^��=��T ;'B������{6*}��!��w*,Z=ワ6}��;�>�=�U�UUF�%�       8  �  <O=6�3J彳_}x|�������#�`��\��}���S��C�, q�VZ�}����_UTT�$�* �y�y��>���z*����ɏ{u/'��^MS�v�G� �@噣�}���{i�ʋ��5#�D�IH�  P     �(P G�K3�9=�s�=�.�� >���=�r��&�J�5S Bͮ��^&OT�B�
UP�P  6�l��9P��ˊ�f��j�=��k֛�כ� ��*��]2��E�.mU�<���Wނ          ���JU#  �  O��J� h     ��*U �i��  #�Ob�I%M     '�JH	S@ h    MQ�1T�L��i�l���@z�S��G�:Hx�O�~g����_Ϳ�gs�X&9�j�9! �I��q�d�$�� �$��$I'�	$��������?���I$�$��2r@$�g�0H@$�/��X?����������B��C�_�G�u3`ٚ�����Q��q`�s�j�Q3m���uh�mWΜ%+	/D�%)t�l�]�y/#�2[�T�B�5rs�X
���)�;p�QM���r9w>�ۂ�ݒ'�%�qp,A�<x�����oP�E^�ZY)MI�x�r�2�;i��n<�4�jJ�<ݛ�n�=���7��ι���s�����>�dǮ�F���)��2B�;�]=r�yb�R�V�K,�]˯mk
���4��Dt'i��{�ᄂnl� CK!��f�)���a�gV߇T���%kw;�e;M:�K��[pU�o�wa�a�&�r�2�~�tt5�}3�{�'iv��W�dڙ�����tWu�P<���
���<�n���b�u� N׎���Vթb8�Ox�T��r�oY;���Ck{Ŋ8�;Fc��^�0���ۊuܳ4Cݬ��#�Ӿ�������Ɩ;x��gwh�C�
!���q)C������TtSf�݃24V��p)oT{^;4d'�����욉�-e@�)j��nn�B��Lo.��o@�%���z}p�d�l��X-�|��Ŝ�vIq�4��7���ǂ86([�=�eާN��׬9���H)Oq ���&p��m:F,�=;�|�O�j��1[f;�6�;{�>R�6^�0�2�ͫ��N�R\��b��"����:*�*�<����`c K8cw�«�;Q��sz*)'u�S3}��^�x.��9�Ɯ㗑ŧ��F��o�.^z�ɝfJ��q�4��x?�N�wy��y��� �{�,��zp����d��n�ĝ�Hŗ�F�3tmE����\x�(�ù�v��nqx.m��E��޻ﻶ �.�]��эmGVn��g%;]d�=8\�s�ܤ��d�cǏ;�ak�u�&��4����,�7��;�'
�|ڮ�
"�05�4�y��.�v>:��{V�'�fHQt]8����͔�0�s�`�(���8G�"�>[/ �kxl�p��.l���x��5e���VF�e���R��^�δ��ݕ�E��\�wEC�b�'���i�zwpu���xH�I��W<c�z���d�ǁ�nZ����{�mW�oݸ"E"�i���42
=!�"�c��`�g5�;��!�&8��&�cm=a�Yz�N^�%���rZ	����'a�x�3Gv"���T�)�0���~i��ĽT�r�h>x�K>���Knj�P�YǸY��!P-Sӧm��.�ѣ���n,�;,F"�-�ۓ�@�;rm�G���!�gv�<2� �K�FY����b����K� ¸��_L�����\Z4ܰ�g�sC�q���Z����#�t��麻S�3�Ղ]S�'�2��{ꑼ�k�������V��0�m>H��E:oA&��awF󉾽��z�i�7u��vw"`n��3w|�!�|2�6�I�2wV1ۋMn[�M�ؤzЎ�x�[�n��I����C�ƪṢ��Vp����Ѫ�[+�;AIs�۽�J��i[�N�(W�r���A�ٶ)�tᙻ�0{��
�L[��!��qo�T\� �q8���6g; 9τ�ϑ�2�L��#�41�ח��^
i�9�'p�F�.�37e��ܭ*�Cܧl��UF�6P��h����a��|{X�ΎWO>�)�����'˄g=�\�5�d��k�w��Ir�!��WjQ[���wx�r��Qz�4��j�۷q�l�Ǵ�K�[@����G����,d�s��˯��}Oo�z�=�`Ȼ!J���W΂^���sT�Ub�0Ӵv�2��Ku�[T�V����Bm[Fmg���jL7��ppw	��d���{�9���gRՒq�B����ĸq�4kCy){��dλ+Ñ:����:Ɠ�=��K�7ww[�Vn+��8E��5��XU�:��o6��qvnn���,s�����)Cw��&�n9�br�u�]6�\���ntsmWGo)�:S��	n�7��62�q�˩$��8�P`I��|�u�M9��OPwFs4>�K�7����d�t�ׇ>��6m���x�sa���$��37S6eT�=��q[!'p�`���G,��w�'](�K�s��0`Ē��e��	l�����,1LS
'����S&�h��hD*9,7��9t��-w�7��iDޣ�3�
4��Wi��"��:�!x�.CwJ�Ԣ� Hy�n��8���N�kzf� ⷬ�х3^��wn�3�7h�7�h{˝�o���gN4���-��zl����4�J`[��v���s���	�)����F�ð���7l���ĕ!���kq�N�Bn���"��8�@!ԈA���,��:]X\j��@wo�.v�9we4q&1�w9ܙ����/�+yh�����t\�R��5�)qۻ
�-գ^R���xD��w(�i�
C�U��K�#5�톋�+Wx7����FI	�V��8���;t�q8Fw]��� �;�H�׍��<��;��r!����s������qI��s�
�$�A��٣��坡�������:D�)6��j]z[�P)�&ݝ��L�ڴ�g$E!2)��`жM[�NW}
ɳZzru=Y��r#���,�M+m��v��dԻ7(t�'~�ݾ��Kƻ���Փ6��p�҆۹B�u�W;ۜ:���{6v#4v�U�Ǜۜ"�:��)9�Տ.A��:W^0��*'�2v[[s��'�h��u,x'K��h�-�M�`��h�A<F�|�x�r�;^%�:�pȮ��`���+�:� D]�������nr�1�6:I.�j�p���m��k�.�zY���]4�rz^Q�)V�d�A1�W���M!G6�y6�������J
nq׭�/Py�A��{�5�b��Ц)�l[�ps�/���Lx�Y\¡��֕����Ǣ���sMݽ%�D#�o/a�e�k���\���aK��=i�T�Zq��e{�����N��侻tm�E���ۆ����8I��K��&9l�K�{�Vc�腅�Qsoϻ���gʝO�������rƱ�v�=2�\g��7���S��uu��'d��.�N���ѨvH����\�M�����&,�'n�)a:��/8�N����´��D�	��X��y�7����D}y�%�	pM�ܐ�*@��m ݔ6�7�O\�y�m�_��ա��owN$��nD�f�S#p�(��3M��3���'���7N�Ǧ��R3���~�M�Q˙��dO{*b�ի�j�z-���C�9��yb)٫�H�sv9-�[�jJ��-K����'4oG޵�Is���gF�٬d·byX]*L��WUbEL�l��n��y�e�9k.yݡr��7�dl��g"�p��	0��KW0� ��]��r���W=m�E5���sU�$�rX�t�	��{�S�16��؀[1g����͜��p��R���L�焤�]x��,�t�J�C�QK�S���l��{qh.]ewhuvr�Jش��;3/Gc��ޯj=�Re1^+9�Y6����y��&u+uC��5Q�35l�f.�79��C���9.]�6P���/A�jw#컷���e�㎤������m�u\�8���A �*ʙ�G�+;��C1���|K�['<�9�T@�֑`�ٴ�03�۠\�[;r`.�բ�����dٸ�gH3vf�]`\�&�nZ����@q" ��ͻVl�.�Xxonk�ol��%6��\Q��٣kN��X��`�g
��ԂB�ZH#�NUFr�6\ѺJcUܮM�.i����]�{��i�8&�)B�9w3�\}u�o`�"��9%���onâ�	����(��ۚ��N-�t�N@@�h��Ȁ��(ɗ�)����;T����y"�s�b�΄��0�YHI���Z�G�\����T��\4wt%���u����$�_ \X�qD���WI	���
r�5rx:�v�Y:l÷^rz.���-y���MQmӼ$[�L}��*��� 7L6Bהּ�f 98n��?N�q�&�D5��9qǷ��κCw�c�V�J�jC���?s ���Wgr�_M���V��]��]a�@8�^����>��罹yt@��$Zy��fԐ-���/�!�b�W��O�=O�K��yv �Ҕ>_D�{q�Ѱ��@�˺Uv�v�y�us'���2f�5�P�$[M���E����:3�V���w��g��;wa�HT/mA�v�������K_aL�Lq"����l]�}�%1uխ�YC�ӤHa�P(d�����z�:�E���Z&�[��5)��"�v��iCuTaz��t�Φ�E��%y��5�,��57l��l	���
�f�[��V��O0u��$��1D=æ)���" ��qt�U�|\\���F�y�����n����s�ۛ>/�Y$�;;y�cxQbьk�$�W��ίpˤ��|^��B;��]P���.�H�)�n�:cԇ���ɣٿj9RҮ�
KU���a��YAKx�j��_)���o�w�M֐���<���Q6T)��h�O8�x��:�h�hn��!�vv3vn�c�I5�K41�N>X�
a<�]����x��!���w�Τ��^N�����g#�A�4�K�h�8t6A����Y֗��OS����l�9�<�YU�ի4>}��H�q��o�Q4�o�W+��e��J�*�u��C������2��ls�8���!�^��27*��z3�T8kձoN\�����6^�XY{E=��%ûy(����FVWFt�4�V�w�:.>hyk��.��v���'����3yt�I��L�x���\���Lz�(�����&ø#b2v��rL(�ӝ�H`�m�)�B�*���/Y��:�\�u,��q��y��rb;��i#1bm!ŀ��z�Qj���p-� �w/bW���C|4Ȅ<��6ӱ�^�Z[�y���^('F�ٸ���N�N�gq�ȇ�wpg�2�\��U��U�v�u�VjsV�	4����b����6a;M�U���悝�ᘧV��ֹ���i���.�z^�p>=�Υ�k˂�`88`h+aBH���	�RR��'�̋�eY"&E�8/t�?lC\|E��U`h���39���7o����v6�y�o�8��5Q�j8T-j�֜����������2N�#S]�n�w���Ӡ>ͬ���\�4ޝ���p㳛�RU�:��.V$�~8ʺSx�T�޹��N(�	���b��P�0c��i�,��gr��	�bM]��yܱSi�8_o$aќ..���ځ7���;)���D�Ȗ.O��ɜ2����_�E�1�C�a߄��;��v�!���s�2�D\������ι�(p1TIsO��vsӇ����YN�����N2x-=ød����Im�m�q˶@u3eY1R���u�gq]&���O`5��鍶�*j�W�	�s��{��*�8�m��d�M��N�cO���y3�� �_݉m������}o(t�X��B���I���"�r��,���&�8��q���&��q���4n�?EÎ�ż���{:<G���4,Z��?P;��*N��bBn�����94	����l6%k~z�Yz�uG���Q�"y��F�YcgeS���P7��$��v��{�VRY�렕�9^�&�{m7GHBW�I�wv�n�;���t�}����1&�1��{v��\Z{���Yq��Zݶ�ɚ�j
ۻC;���|�wq��Wd��Ũ[���@���(�h�:�M�@H�/����}�K�&�(/_���wA�>8S���n���5}�]���tC���k�[Wr�8���!v�����V</�!�8�~�#P�̭���7e�\=�I�1%�1(AjT^EE͘;����V�r�<ʇ���f,v&���0��wA�w���Y�y��j�Z������K���w\�´�̹�� D�r��no0@iӮݒd�EOi�ԉ�tYw&�L|���b�]�˳�p4�6�� 50�hٜypES���ήC���S����r�`>�ɷK ��2�a]����I�4���Y븱��P\���Pu�*��M�q<5��M�tQ�g�]�L�ƦNs<f��R`&$�.T�{�畟�~�օ��*�\�k���fϖ�e�6��X!� 
I2���v����/8�	�E��r�'�p�G}�k�RQ���Rop����g|�Es���bqG����'��G4�k�p-����' �L?�(��٥׬[�T�I8��.�����(�[�j�3�D�	,�*���.ɕ��[8��#D�W=�^���)�p���F��N&D�.!� �������C{�\�4r����G�(7��o��;�q�פ.='����:��@ǔ#�x��	໼���H����q�o�ĭ,�oP�l؇N<G%Fv��q��ځE���>�$��M���)��y��M�ڡ���s7[9G�b��L�)��f���v�Bʵ&ˇ8�=�u���V}��I!�Y��!N��;6Eòc��:�|w�y�b��pw�;a�&E��a}�7r��ӹ�e��s�f���ecF�n��n]�+�R��D�p�ɭٷ��;�;��i�����M�wt��n e�Au��s�h��S�&�A���������2_�<��Ek��-G.$�M1X0̺��j��o?C>�ß�^����sh��u��c�/6�X���=,[����z}'��N�u��[�׮1��ux��ۉ�l�S
k���:��-��jC�mt�ݤ���m�p�y4q��6��};u�v��v�GNl�+�g�#n͇�=A��D���9s��=t{���[�N����?&7`�]�d쇑�۶�v�=�t�=�1g7N��څ${��]��ϫ��AɃ���kc�%�=�6֛�Yz�׭7ͷNB�lgOR��7^�hڌ���Е�t�j��xz�l��ms-v�9��9�a���l���	ý�m�vf�2u+�G�oN_&�;gTn��o!d|v|ڎ��vN!���M�\�#ngoM�K�^e�V�q�U��6ܼ�C���p��;[)log���Ծ���d":�ڙ�.�Ij��n���q���=v���n�ֳ1rvm-�����n��%B;��8-��i���vw>^i ��1K����4:6�l�al���Q�϶�]bö�J񋜶5:�u�^�� ��]�!��ʆʖ�t��ALR����1A�.���rm��vH��W/���.W`V۬'n-�c�F��vpzݻM'%�۔g?�?��������mp��كe%��)�۶1k5���)��֛�HU��s�5����v,t�D��D]˶:�łA�<6��o[��P٬��X/D�bvl���'Mu�9� ��ݺ2�Ct�I�΄��F�ZŃ���ۓ��K�H�O>����K��z�A�%{p/F�ucj���$�Y�@�.zk<�=YG���˼����d֒�	9�Iܧs�e���H� ��o�/n��w�1��K���zK�%K���Kzy��ƅfۮ1��la�E���=cfON�]
�nN��u6M�=oh�4���룓n�tW�vv��C��F�G����guօ��v�b'����;/}��u������	ԩ���\�u�0�^;Kr�9�h&�6�M�.|����b����;��]&��=����;�h��e�g�st��+�*�mxq�abHng�ғ�`y��"��ESJUs���ꬵ��g�����Xd��G.��?dpʜl�[vw2�֎�Y�l�P�,�C��8st"Z�����n�f�v�nּ�	�R��˔���㫝�;P"n;n���E[1�Ϯ�͞x��d����\�5�le�������,����<�.�m!͵�i�Wt�^w��s��{��t!�髆g��.Ig���R��M[]��g��v϶l��%6�ۥ��ʜ���lm-�IV׷r�[�p9�복�D�V[��aٍ�ݝ��wce�f㫗oV�;1vzvŭ�]��mtf���:���;c;�Z��.�}��]�vN�8,q�gm��=7�`����WÓ�rwn�h���
��έ;qr��F�Z�6v��܃�F�F���GC�m���n�NѲu��Ϋ�����udM۶�%����b-����]l�q�nxS/ph9m2�r��t���ȑ��ݢ0�y���{k��h����cs䭙Xۧ�Y���ܾ���4������۷mmoBz��%%]��ۡ;[��ikݔ��{����n1�F�d��#����gs����&W^���άG$���C�ݕ��Kv����ۣ�N�$�<��p��r�5�z�}nl�ui��g�C.�n�W�n�m��ہl��t��F�X6�y̯C.�z���|����E��=p��J��7n�����Gn�j(�1�v�Ӹw�}y�o���Wg�{��l�{�<h�z�&ƐN���[�y��<�ەS��vݸz�y�X�{[�ǅ�ݔ��^dw]ng�K��8s��lA[����K���`��f,�Q'|��`��y��.Gr�����fu�ml���{A׺�����c3'��{V�[�զIϫ�[�x�u��]��0�!�۟FGgUtcq�+s�u]�y���u@tOmI�-o2�悖{WL]m1<��/CrB���%����`�F�n;S��X���)u��f�2��ݷ�^��IZ�*���m�j���bK��^7&ze�bk��1��^��4��v�t�m�<Ɠr�q�؞a�.�u�ɭۮ|G��l뉳���1�m����.ۨ�lfp^^�׷z�Zf�<���c�uJ���9C�u�ح���;��=��v������vz�Z,/��tk,��[I뇊.��bxs�u�������m��N���1�g�����/�<j��b����y!��]�4���S���;�-�{w!����3A�d��żJv�(�/���V+ܻ��m�c&ݓh��^lX�n˭�V�ۮ������.	�d�<q��.�2pܤv��w!o��'!��Li�n��y0�����N�v����u¸Ϋ&���%�Cp�)G�1�����ۓ{M������uqUu�u�('5��<f:�ŷ<h��n�l�ٹz�j����w<]{`�^9�NS�ݸ�u�J\POA�ˍ����k��sQ�5s�|�=�k]׺�;�˛�� ��X&��%��q��E�''��^{�/M��[���O=��N:�n������6�#9a�,�G��t��ڲ=��M�#�c�k������lZ{k�!���χٷf�-�'Gn�]��|���3�y�ܶ*k=Q��S�F:��+�����v��i�Q������ۀ�q��}�r�˶�-���k���s�f۰�<8Z�Y��۳G�i�=�`��緇=W��p��^r=)\f��j[��17s�]([\�֜�'�$e;NS\������v��m�����t�����q���d��ۻuNQ^/<�d���!��
��/*e%����$4��wa�ٗA�f$9�����<�/fN��9Y.zh��TQ���m�nݮ3�yn�ag,��ۺƜs�6�#<7<�7���X�ll�
�8x�4u�uW �Yܝ�q��v�2�c��s��j�df�N�9��ns�a���n�����\ވ.;p���v���n�ő�կ�G��	�*�;���X�mk=\g���mgN�������nBt�p'8�'k��C��']fl��,����J����vGm��sr|�gw̆��ҫ�:Ih{U�˶6ی�O�r\���y��틎���\p���;*7$�g۝e.=r�<��ؙ�i٩7H��;t,�L����=\��lT��f��=�ثo=gh�k;�����ճX.��õ����ڍ�q�%�NᄜG[�������N8;O�Fcx��u��i$�S�z:nv9�ի����$k�yᰌY��nu�;`�ɑ����5]��wm��#����q�s�74TwH��ٻ�{	p����|���7G>�a�R�&�m����k�w6�#�]g��	��H�O��;uZ�PV�0�d�l�Ȝnx��Wg'��B8.\vѷZc��۩�������]��M�*t��lv�^.�)�!�s��,��<��07do=��]E�ѥK�c����&2�q��m+�u�k�����k��v���u=�����8��6�ў�Z�7k�Wm��Γh|p���9�v�:�[j�v����瓛v��z�ųr��sl䴅�;�/g-�!����Ѭ��.���x9���>�oϺ�3ہ��u/Mg���b.\47�z�㱷��y�9���/7��c9��Sm�<���;y����>rx���6�81%���-�[��,��^��X�Z��;ю��v��rH�`ٸz�ė&j��:���~;}��M�M��̽�'d����[�d-�vζ��;������iܝ����ܶ.c����љ��.׵֨�G=`ѫ��糎c���VAl�m�Uu�I�Ým�U�紐[�����X�]۵��b[z87�=���6��c��^�OVB�;�Y�G\�O/C�k��zsd���6��j��9U�68�qq���1ck������k^�f�ό SA�W���g[�gM��5�a�l�`����vRɏ��[�@�Vم���a�Ś�Sz�;[v�$���=��\%�zu����uf��X�'\�91��.G�m����z�_S�S��-����݅�#�u\g�������M�9ȼM�v��4V�+����T�,�&��{n"��۬n�5�`��	��v��6�n8���.c��+G�������g*������0�I��g$<V�k�m���V!ܱ����{.^����yקlN;g���;x�=�]�����lp�NL�狇[��'A�*�쥜��s����K������M�V��|�v��Fcۄݝp��RUu��;of��\[۞4��~��<{hՆ���,W�CL�-�%Z$[n��m��}ﾷ7Y��B����	��Y��!9<\�-v��6;m	s�S���N����ڋf+�;p���n��d��D�1��kc��l%/j�b�tQv,���[t/=rx��q�u88�=�����t�<.��!f�8���qv��}���f�km�9���뛧Fvwk��UiVqt�+�A�;N+�k0[sAd�ٸ�ݮl��}�}G%�n�9��[5h��݂�^��[XF��"Y�v�������i�ܺ*p�ݼx����FwZ��v�Mgl�:����3�]5v�l��ǬD�Y��d�\�@>lq�d��;��������-[�4qwl����l��JtH��"����m�`#�Mnq��\n�m�ܜv.6msئb�v]ڀ��}Ң�ܘ��!n3�*���)�Sc���\��簐R֓ax{]v��k�����]յ	:Z4�����n��9��To����r��I�!F�U���@�8���]�\3�Ӳ��7U�c�V�Ù�v��N��鶔^�K\��	�a�*�a�t5m���9�,\��z�z��X˲X\-�a���ΨԀ���7[BBѳ�Ӵ]����v�.��<&��[g�;[u��-�7����`��ŊƬt�;r����V{T�F��Эmۢx�3�7`��J�6�{dy��A���ST�V�z��%.�����:~q�x��n�Q�f��'n.���������'� @�I�����'����|�c����۬=!��s���y�4o�gb�)��2X����d{�;/f�������X����ԝ<�)�j�
7E#4���s�����9��n�E�9�v_G��v`��*�{�P<�3q���/������bKsZ�����-�IjL�ӦU�tnaN�H��a���������Z�o�Ⱥ�5��kx�J)���ȓ�
�1��^�=3���h�>�=�l�=5����1N<7�f�l��Ze ܺ$e#C_�Ť�MUn]��������Z����cs�e���H���E�F:3�6�o����IwF ���+�8��/{Ô��`��1���bl��Etu3�SSv�c-x�p��N��9�������y��ؽ�����p��O����$����Y�Ma�/a��V`�S�X7�+�����Ut�|e��P�ä1��5�۩�{޾������ypq{$\��5�w�)"�"%�'��x���q���w���;N�x�5�R����������/˜���o�K��}�{��.��t��I���m��]L��d�`S�z@~6g;�����y~�:g��7뾸{���e����0�}��Y��=�����ސ��p>��T{܁�P�����b&V˪s�=���t�}���`�H���ՠ�����}'������:p�@�n�o�r�p=�'y�|W��g�.�q�3~�9|k`���p;
�5�=7������t��.ڳ��gCd�ew���쐕��v��>{O=C���9�7�H]u?y�2f��p���Bn�������އ�x餸��|�۞]�K�e�z{=�Wx�EY��s���z�햎V�-_�q�w����?[���4f���C�jՌ�f�'wx�^��wV����T�N�nf�mcׁ1���d���໔�tz�����v�ЖOr�������8����姫��:�= N�u;�P�'^���*�=�w^>�D원����/���Y�/+�ϳk�u��^ ?j���N�Қ��Ic37Bƶ�B��ĕ��Õ�ڴ�ଌ�F��t�[�Eنf��F���s�u�;�$K�F国��n�α㇮/z�ק7��>�i�A/ګ�Y؝��D�3���?���5m��*ӳ5�P;��E'�>ܻ���������d��L��X�E���,�4C���W�b+�J�{��ʝ_5�zG{L���w������\��U�<��J��D=��4�P�⛳�!��va��/)�v[F�OF��mk�ў��Y�W��b���{��g��pǾ�w�|n�.�3����$/{�bU�]�G����-S�o�z!�ID���כi���vp6��J5�ʳ�hyc`�w�����/b��oj�Q�r�\������t�|;}�b����}���7dk�g�Kz\��z}�^8�T���ƽ�ı[�y��En�c6��\dU�G�7���t��&���|}c��n-αvmcU�����u��S�bW�槧��w��>��yg#�;����`����Z�nJ�>ه�ٴ�}��Ak���6��6����/���PU�]��'���`�h� ���k��@�%6��Z�q��n�����C�7�q�XO6�L͌zV1V+V��u�/b�1�`�%��w��X�RR+-�N������66s|^V`�՜��⛞��@�N�S6��{�������7ޚ�|R��h��-�Pnu�OZp�T��GF��W9e��@�@3�7ܽ�qfٲ��Ë����>��==`�q�f�������=t-��ӯm����ٯ���a�r�-}k���p\93ͱ܁Da9�B����d�;<;e��娏�X��7O��� .�{'gJ�<�0N!,'ަenv����ʄ3k���E�os\�f�����fﯟ�1��Ðz�1:��sه�g\���}d��W'+q��c��b	�b��qgH�'�Ul^�Z1 /�&�1QR!�R]��즈�x����o�=QHx�i׋]�E6&sZ�mq9�.0e���͘�,����0��x8<gS���;~��`Ѻ�u-�l¾���������S�v��7@�~�n��c�dQ4��!�x��2m�wrT�k9A��77;��{��,�g��N-�	 R��k����Q�/�h����Y���ct��N|OG�'���>#���ěV��NJ�y��;��љ�P{(�X��0�T��g'�!z��h�39�٦}�{׸�qꞥ뽻<�Э��y��x�lD�;�F@�5���>���Ś��sۍ�P�����\KN�����4{.��
��3F,�`�u��7D�q��nE����PO�_X,-�{������U4H����;�si����� `F-�Tc�w���'���Y��sض�!���ozt��%xx��;�:�.`yI���ng�rMz��P��{,�/������o����G|%~8H#4�Y^���{y0c�Źp��7�8��&��}���n�)���=��_^�I%���{�P\�<���9�ٔyo<����^�^�M@���ڦ��D�)w����\_�=�k�û�%��3�8��C�5[1�� U�F�1�J4z�-�$����9�>�z
ch�[;{l�U�����y�;�i���������	M�w�ݷ���wi�n�O%'��8��בD��n���d�Y8x���{_� Գe>yN���HJ}n�l�<(d� ���I7QDMiXw��6>�����G�W7�)��a��ctaӳ���0Px���<�����R%=���8V����J�E�%��o+)�0�g��@���R��5�&��)�ѭ��g�䋃/�Pa�n6wSF�f,�'�e񶞛g�pҽ�9�9��v�Ȃ����#�%=Ɂ?^��F\�fpԤ����-}����F�:���w^I5�|��t~�>wXt�Zz�,�W��m�7�^-e�����s���F\������>j��S��|��N�^5
=�|��x���J�� �;��kۯ}K'��Ɓr�a���:5h�=�s���3�>�p�\�L���f��ބz��
vi�4��W�ѷwx������qd�s{`�;��	�f�����|=ؐپ�y��>^>��z %�;2J�ם*,MʁJv�f��m�D?lT<t���aPDcX�^����ȡ����;���_a��n�)�xzYs�K�VV
Ȓk*���*J��{�q����$�sV����uq���=l2b��{�[{��7c��Ox{؋~�t[����S�[��3�	���|o���$�pi�a�sH�ݻ�|�m��)���aO���f��9��K��t"w_ox�\���o�V�rf��t�!��<��v�����m�{���v6�{k3JPN�{6�oL⪜��rպ:��sϮ��E�n{._);NG�f�Y�nm�U��f-���3/ظ��{+~O7�&��޹=k����eo������Q�N-�7+^n�-f�8C ��ë7i�Cy`��d\�����g��]�|����齽���<�_Y�^��	��4?w�z�vW��:����v�߽e+ld�~��V��E�?<օ]e��ǆ�0H�se;�{JS�os6UV���\ƨV������ �+�N�yr�!��'���\'��Z�����F��F�����guC7��Cӡ�YȻP�9����w+��޵����]�,7;�K�H{\϶�̑}s��k���=��;S��>)�^�^:^N������Y��i]���wrd���L�����!��ۨ3�z�L�;ܝ�+�PY7�p`�7�af\���;�}�(غx3����p���7��z� ��ˆ��w���+�/���vx��gH1{��v]9�oA���p�����7)��������ipja���C��f')��5�L�轠�GXQ"�=������^�w�N｢ ��^��x�Q�#w�/�S�)�z.&+����gwu�!��b'�gws��-���9�u�}�+=�����^�]^��@H���Ni�:�9:�S�P��g]ӛtّ0u�R�8ֻ66l�8��p��+ъ�1Kˮ��Q�9<�u��^�g�����hX{rA�v�U����ɹٻ��9����[�(?��)m2n\�:r�=�Jɮ���%���H����ה@�ca��^���f�21��vy��MwvLO����������ܚ�͇��{;ɥ/x,���ʂ0mggX�1�e=���	N�ᛑ}��܈n��=H�:͞� ɪ4ݘ�ƴ��x�h���V��*��Y��'>������M�Ӊ�i��.w�|(����۵�e-��ogd3zp�!3p��VP�~2�.^~�����o{���%Qp\�_���P"掯���2���Ӊ��L\�eډ[�v�W1:�<I��6���z������}ر�F
�7�^WM����y���.�Iߑ:9��۷���]�9���y2ϳ�˛ }������:�6똺gJ�M�qz.��z��e:�o[�qS4��F
��[�|/�U����3ȮO֛��:x��~<+��.z]���z��%��~�S� h�G�ޯ O<w6S�O��DG����%��ˆ�������n��yH��v�b��VCy��������ڼ1,�{��u�ao��c�������K�s�j� ����,�u���膔��S}���>�J�lg _���{��9e��}�'U�w�r�&�K���Tw�q7��/t�v-����,�??Z&�on��ݹ��7Q��G �Ó턖&mƟSn��I����F�������<��	:V��`�Ԝ�;����b����P{��m�m��Cle�T���NЇ����v4�00b¡�ˬ.�S�$μoJԮ�hp�E:��[Fa�`\��ꍐͼb�.j~k�5���ݣ���`��p��`q�&��Wt����i��d9�5��v��!�3�>)����gd� ��e��P�4a��Cڭh�1�����Z��֪w�ʷ��n��Pf����(2yS.>�祐�<��)�m�%�O6ݻ�H���{8�Sx��<|G��@v�Kξa׃s|���١nN�]��̿n�WQ����a}��z&�R����>��=ϑ���f���� <cSC�{�g��9����0��.�
�q�|��S�tvG���5���po62���(�z��$b�F�̈́����C[�����jv�/x�����;�õoX��=�+�L�x��R��p�N�03�u�L�'��˳�������u� �i��MI�f2�����4w\Nbʱ�J��``��pF�VIv�(k�{Ƿ��޾ٳ$�fkm^Z�qd���u��Y�7]�Z��~\���[�e��L%s'ܭ��u�3�3y��y=�r�KLT��o�csJ9��i3���y���%���Vú��sC�
�x�\7��S��%6����,K�N� �4w����&��%N�:+tv�ܼ����3�ٽ�|���Y�B%)�u��b��El��&ė�{q��BaStd��JcB~�k�
�AN	�����HƗ#;le�ILe\II�Ⱥ�OX���X�`�/@D>Z�#8�I��n�Y��e�=.��wL:�{�T���+u�v<W�DfG����U��ֆ�t�y��Yk� �j��>��>�s�㈋�'zl���MN���d��X�|k�t����r˫�g����tM'�<sX d�E/m`a��Ȇ�Q���7U-�.�K$ B����%.<�lw�M]���gY���	)�ok���Om(�iH�懦ze� �ї49���ӯ�8��<X��O��C$�=�	A(y\�a�<w<�s���sU������O$3ېw��-^M��'bS�t^<wUHG;�x����OA;6��_`��l4z�\a�����^q����Hga<k���y��0s}��MlN}F��?jY�n[ � ]w/�mf�٨�(�#ݙ����n��۠R:{��˲abWc�~@��<K��Sw�Y��W���UP�n=Ű^��We�ˊ�����J;9�y�x���<��"�vj�윁����;7]9:�^���Y�Ogs�y=:A�=d�mv��x{OG��ڼ��rï����61�rX���4�+���7hh8ߺ��3�ա�8.��K�f��c �����n�%f����M[�Ѽ�3�(3.����7�x�_�����|4�zx��n���Ƕ�<�l�]��8�n�ڮ@��9���y`]J�����x�5�u~�6觏������eצ
{ux���T�������Ȧ��jm��f,� �ˌ���5���k�v�k���8�`�fve<pȱ����'4���F
Ŧ2��t0��d�N0��pI�|`A��Pñ	=��E�-fLdߚ�`�v�`�0.�mv�7��������j�}�5S�B����q��˯R�Z�j����:�ӺZ��Ѷ.�5^}׸�W�!fw�����r�J�+ct�9F��7VA�;���h�����p�a���E����b�g$U��{܇{e:����3�=���8�2��=���Tp0�d��e0"de^�[�*�5�ӫI�1yB���:ν�4���g���U�ܙpE�q���r9V�x�.웯`��+v�/=����
����r�	�\h
{nWo��8*��B>�t\p���4 ���<��������G�Ü���7�7-8�\W�d��󝼭�Dv�oMKQh'�ύ��T�$�N-~�=�����Q���wr
{:�3�L�Y�p��5�2�&V�;.epA/��Cx[v/g�ȳ�p�Z	j^��=�Խ�2;���cq/?t`�<2�J-胨c�ŭ��əi�˹����&�-9�a����h�����Wr�7vY���K��G�_I���ޙ��������b;�jk��M[�
�4z>��H��d��Q��R2'�@�H��7#����\�wZUڧ�b{���jY���:Ż�6�K���;}��L�]S���\���^�z_*����ziʣ���Y�Pq��!�[L!�#��o+�}����e��P�7��;��p�/w�Q2���}3}N�|WgY��@r�G�|�U�I�����! �I����k�O����}��_�;����_�gBn��V�����$�cu�w;�q����qvz�:;V�]�U���2u��snݻ�}լm�޻Tdt����f�]�Nv��I4�im��3®�+n�4Tn�^�q�pO�L�|�'�<�Wm�;[s��x�'��4
��`�X�d���]����&(�l���.�f���r���%v���ݝ�I��'�3���q�ӛn��j4�9��:�uQˍ�@�U��&7^�&ݺ�wFP�O�簻��̗.��ú���ϦZ�)��[Y�1��;���wBvǂ�v{��۶���=�8���ۘ�����[<�\s����.�5�ͮ���r�ؓ�@�n�=���9&-��(:�MȏEWx�p�ɸ�5M�ڬv�������n����ex��q�b��7佑��^�gk��D�۟@�r���ᙻU��=^;��i��x��4��L��<�m�C�%\�z�`�άm�J7�6��4�<Y�=������-��^�m�Ps�tm�w�u8wm��y���;�F���:���\:z\��� �n��)�.9�m�G6�K��z��ŷ� ��sZ�kf�\v;\��q�8ڶi�����v-���0J�,���.a,[�Ƹv�;p;������,����n�mhyp{%�]��g/B�6�=m�c�����0�kβ۷��]6�ˢ���k;gʸ���=/�rcv+���	��=�捏9���l���{7Ǯ��!�(�u�ϱ�s��qE��&���&�"��tQ�j�yl����j�f����-�M�X.ݼ��LZ�rs�*���6�ùEwk�v�CGn��g]Χ�S��]������n1�3Vڭ�k9Cx{�C�ی�[<86��a}�+�ܗ�Wh[<p�m��`�.9��-Ҏ�^zn�0[��I�۳��;��v�9+�Ů:N3�kn�o�s�6˰;��ky��V����7%�d�\��\v���*�
�p��ٝ�Wj.��]Y1�_X��6��e�غ�Ħ{0�&c4�0�Pҳ��5��3�Ι��n�ᢲ��� ����խ��f�7wnpէ9{�?h��k�w(���`�1��j��2e��>c�34w9f�y�>/Ӛ�h篩�����ѣ����^��H{�wKQg\�2�g�gM��Y~�J�;s�w�r=9�t⽾?�C�t�3�����=�(M��ܘ>�"��ǎ�J�]k�wA�Cb�2�-��N�e?2p�&F�Χ��` ��8=y�ޘ��B��\�:�k��3�MY���u���N���QP��̙euk���h	{	��3m
���7�笋��fݛ��Hh��ٶ臼*��\I�2�;�a���"p<�C{��B_l9�G�{;{��l!#���:�)��	|�3�����{�����8MI��~@iA#�ftiW��<�b����t���r��$p�&�IޥMOP���F�8�$֪>�y-M������Z�}=6�©��7�f�b���㫶�c�z��l#�
;r\��{���D���Ď�[��ƻ{��d��%����kvv�\����s�<��T_���ʧ��0�m��/S�dҨ{�aY�����T8^7Ǒ<5o;�m��=p�I�S�5����D�t!r<V�������d�x�:�tsO�.�&E}�IP'^Ͱ>��ʅE]g.uw92�{���p��|�	���.2t���]8݃���r-������ Y%��:�t[׋i��q0��3��dw<��d1�jT�<׷�v����M�������O��<�۬Q�va`y�d1��f�i�i�=��Og�N�;���/k���M�۫.��n�]�0�n��۲ez����99����^��@wb[�'/`���`z�����w��{mݬ�9�suٍH�::�>H7\v��!��q���y����#hN���o.k���.��ur��i
� �T��XU�8KN�d6�����ܜ����v�rpn��N{oc��x�\�(w�$o7��Z�1Z7r�|��P�[��N��F^�1�Sa�p,a��٭W�F�o���m�tm�||�n��~��RI�am��p���Gvl/�9O/$S�E�32�g3Z�|���_�
'���A�_}��~���������UG2g*������:�p��c��I� ��b���ڨ@~��{6|��To�5���g �Ê��@�RF�*H�!���v�@whZ��:��+���s՞j�zl/0M�6q����T�]aw�g�pY3-O���pw�B�ɍE�>�X�� PIf��:w;4d��XF	��erțoLɺ��%�O�\��9��&�
���Q�5�n6��;�c.5ϫDŽ麇�S�������D�UZ�޿�~2��q�7u��H����ۦ�.�ssu�vQT�0�+@E`������w���R>�H��}�M��2���`2&i �VV��Ȥe��c�6w�߷]~/&���9�e��c@$Zٻ�Er��-t֋�h���^Ǣ*�h�20�gF�x�&�)"Kj�^�����F���fҳ��K���n�DD>;����X۲�;u�L:9�/����䭍9�f�us� y�����3�u��.#����uiJ�j��X{��]e=3Z���<�a���q`��N>[��B����f�t�U��Pi���q��Y.BP�HF��Q޵�2�L>��뻷�������������]L9��H�8�`�[�a��-��خtK�=��;w��{���ы�D�U�\u񿅜z�-�_o�����DB �D.�u��:�wr"1$t�$������^� M$)�`�˻Y}\{{�puZvK`���*��}���Z�]�ⶶ^����([��dw��r&��0��1�+ً��%����s�ku5,�N+n�@���L��I��F��m�hN�F��O][�ݶ�0b�M3�yuhk[t�Ke��'���ų[/�E#/Y�Gx�WPݽ�����	�2�O��!�LJ(#��qQ���l�UE�pn�2�d��vɼZ��l0�ɳZ�����Z�QP(�ւ�4�Y�.��?BS\��$PH[Pb��	;�׻��i���b���~�o���E����b�F�9 f���D�9wP�0���LM3,����="�<gc�j�U�ۮ��N���6�1���3����p�b�h�9�u���o6�A�듔!����A1�a&8C�}x���kﻫ(������^2�ާ��� ]����λ��ǎ�pP��G�S�Y��8��xz�+����yx��Y㞃��A�]�)F�q��p$$�d�4BŽ�y�J�^A��C1��9k�|�lH8�)H$��y��tG�/F��8S5DkU�Aχx5Q�*(�$�2?�v@���9?ffU�^����d1]��C��0�$,��31�TC��q]F}�����Eߡ/�-��H2a�*�����s>�;�տ�.Ht�W�^H�k���ݸ�g3r#�YS��r�Dٚ����r!j�{�A_U�~a��Qv9���2T1c/y��0�v7���M�0~S"�U��a���#pدV�x�M��Xa(��7;��N�[�Q�x�ٽ�I�:#s�Z���Z���:�ۀ]��ͅ�ǁ����a�H����dli2���njѥ�v7m�lc�u��nÚ3�:]�%�{/K��.�jسX�}��m瞔0ܬ�y��ܐ��;x����[b��;.�Y��c��֞#$�簾ڮ�qݸ�`���Wv�yKw�|y�ɧu�wp��3��ܪ��F6�-r��أ�E��ϩ{���/���u��l�$	ʘ�i�]�8Ӻݦ�,[
u$Zą�q�`�Hэ�T8�=�un�C�h����e�[&�Ri�r��l��{xp<�[�<��v�.�{�߭�Ϧ��.��e�� �m)]ÎVc����<�^Fe���m��B �R`#�P�}�y>��.�/ֺ�F�vfd�{�˦���<M� p��2V'�x�f<� p�V�t-�o��ʢ���>�z~^/
�qn��;���a�`�>��)�Lv���nlk��.v/F��&v�ִ��׿_���kv��ì��*}�2�f�\�W���kR�$�D��K1(��	��F'�م���QΟm����U�Qyы�r�S�R��cq@�o��v�)�S9yW5�m��!�H���H����tk�����&��8k��0r8E�P�@�ض��gY�̙6�D��L�f��$�6P���l�~*}
�ٸ�;�{+�fe�r�E&1�La!H��$8��9�r��߬Cj�]�s��3�~^�U�x��&�a��m$����n�.���Da�S��"�#=�2mU|80�u�0H�
&D���r=���o[�W��6=a��9��s�0�q�E@�2T��Ée.���kdתM+f�ٶ_xp<����h8B@h�
պϣ�ٙ��o�E�1�bG�>�ʠ3g:��� b8�iƊR�<�u�]�@�.�ӄ�Ô��c��e��3]a���äu�"�3��=׉����y�y3b�<:���{-��Yt���ٷ"�%�K�o9\z,DX�K.�͸���wW+����#H�i� ����c̋��sG>҂��,�P�E����@o:��f�G�r��ٯT�Ǣj��6��Ѩ<,�J��m$++z�������j��/ֺ�F�[Y�����Y�n^�XΉ��0�ɶ;g�pm�u���st.��5�W���P�[m���^l���~���Rj�TM�b��DFbL�5DF�z$C�1�CH�]f�>��}��H�I=�R�.yl\��+8V�`���$@�ŧ��	��xa��e����G܅��XY鋊X�E�����羅��:���~�e�!SM��mt�#2�oݢ��j�^]���x������]�:m��펻9�
��:ô4�fjI��n�vf��S��=�H)̺ŽY���:>�we�:��#��p��b��]���g]���5G�鷗����l�d��c����F!��ٙ������b���g������^��+�Y	% �[���m���4��F����usՆ�k�ԁ��^���[�^�~S!�-��ʴ�������M���$Y!����#+1k����{F����=Ƣ��" ����I�_�M����Ȣ���{�+�f������/	m�Hٌ��4��b<��g�Y�54A�����f�EQ,����V62B��6i��	�P�ѕ	͛&q���j͇����mK ��M�susb���9k�dOA.uWsZF�ʞ�7G\䛉�mPkͷ��{.ɜ�l �GEܙ�.[�{~o��z繊�ɮ+n�K���|���ۧ���
p�o'����������.5r�;�M����'s=`�;m�|n7v��Nڲ�ٯڶ\�9+�[�A3���n®z��uc�쑫���=���M���s��t�X,����L;��b4n�ݣ�sk��A��pG=<`�cXs�8�kk����?N��	67a�0ԥ؂촓L���j�A�&��*p��L���4Ou�� �BHQ4HD,�I�V�2 ��9�]�ݠ�&O�o��5<ez^�1��@�E�v4���N���d��n���������*���32����E��b8C��(KL�<moݙ� ͜]��L}�j�{��<���|��t�H8!F20�k����"�Gb=k(�,դq�ʳ��fFR���ܬ��;ك����+*��"��>{=1v~�&�0BL%a]cǱ���|Q�ܛz��ܬ���bվ����4Ȏ�2��2s�nxeq�p��/[��v�.�NJΝ.�N�"<,�J��m$-���d�g���dW�{֭b!�4Z�P��J|LL�n���\^���W@t�ٯ$*�L�<�ܬ��j���Oh94�^Z�uV�w��ڨ�(L�𕺝K���ʎ7�)��x��(���P\p�Y*�f�0��}��_~�ΰ����H�I�t9w]���s}���]D� �IIQ$�����>�ǌ��x^?�,_j����j�I(�c�LרѴF�1�]OI˳��~�d3�Xc�E$1���c΁\�o������Ȣ���{���1~� ��Y����&Y���7vz#�{�ذ�A�6A���/;
��. �@Ќ6�v��s��ֈ��v��m����q=<�.��)%����,co5j���b�s�֏��C&N)�����:��B3m5jθ;q}��N���7Vvz��M+�C7d��&T&8��x�Gf�+7Y����-�Q�q�*�Qť��W�3��.�b���i���'ݕ[:��`�d́�Y �o���;E�X=爝�>�+���P3�G���� K��N��:0��}�^R�ׁLfG����/ �·7���|�4�PSr��n�gEQ��d��Z奨��*�,�COo��p��,j͛c{��쵘 ������Zؑ��i�]v3g[��70�$��G&j�@T3酻{�i���5A��NC~���w�#�LR�gK���յa���y����	m�\���Uf�qn��-O�����ڞ��A���rԭ�Z]4�
G�'/�ö�}��Hy^{Έ!��"��Y�6��ݫzQ������.����U��P�OzQƅi�+���Ϯ	g�rTn���e���9�U56!�u�|u-Q+;�RfңGig=�� �]�UO$��eo��kN{�fK~�/߯_H�"�B���sO�L���E9��{=�À`]w}�B�b�������zȢ�Ǡ����vh�N�[�R齅�<	3)����P�n��u�����vq��Zvicڜ��Y�g��g�"����;2zxגi��W�8l=E;������zmמ�YU�~�k{
�p&0�y��Y�\��>bN�j^�]{@��XS�S�Ld�*X{���ø���!�/��'�o1���c�C}���V�n�oEf��Ycj�ü#�@/ /��I��7��ѹS�&m���~��(��K1n������ʏ�Z.�z�U�91UI��W5�(�{J:�E���Y�����P�O%����<
^^#S�Pyz
����9a���M�x���Kh7�Tś.��ķ�m7Y��E��Y7Q�Ive�P�q2�W����g+���^���w/gs8��� áhy������`Z�lȤ�sU".�M�%����ƫ� �J�L��&pB�IlÙn��j�'B��X}Î<�J(���B�YR�7�l� ��}Ѧ���xH��v��nU��=<o2���9{O�7[��M�^�͓�Z�
2q��Ky�"����N��\qQ�9�y�)�+t�v���4��+ȍ���Ҿ��ռzC)g��A~���>�]g6/I��i���Eͧqe�<��X�����i���`,����Nص�{:�JeA�ba3lo��-S����k�ʗ�r�Ǽ� ���-���g�ps�l����];��㦟[]/�E.(����5��sϺnP��R��{��e�ԃ�3��݌�]H�
�vG�C�ˏ=�ٻ��ɤ*��$bK������ͭx�W4����2v��h[��]Ϟi.y��wo����}��ypo���V-��P����{�0{rI�6=���t�iW�p��w̬�}�4,;�f�U��x��b���2Z�KZ�����r5�캚0b��ʹ=�ۍ�7u�J���%��섆'u��.�,ĮX��PJ����뻜��(�Rw#$8�Cy�[Ͳ�hR}»��H�>6k�Ӟ��.F�I
E�!����� i;~���i)_׊4̦���ՍJ�Jf��Il�W�Q��j������E��JG֓L�S1�h{�6�u�B{��������y�F��}�XD5�B=B���G�ƶ{m�3� �f��]��[�8�7#�Ph��m�O6�p�a��v6O��z�cE������#��*VmϔD�����e��C��>Mc����l��t�A~�H�qI�u�CZb��u�����|�N�۩��i)�_oi����9�v�ݪP����d
���TX�N�<�g�X<Y~ UU|o����>��=���v#�(AM@��
*n��
�(<�bՙ9�r���>�[�)uZ]v���Z�o.�#|����*㷩۷i�ə�p]�oN:����d��:YP_>�iPW��+}чhUmi����C��H�c��� �|D� �]�sAhw^i�2����D���U�ϗ_׻;�1�b�!Q�pC�2s���vl��@ '��A�#�!��J�!�2}��*��0CH�q�ڄ̀���!��ݢ6�ې���v�ħb�8��Ew������j�0�&  ���uE)�4���g+����Ug����~�~���'|TG
(�a��M��^I��g������V�ς��w2�ķ> *��3�<��D��Q0ae4���e,���!G� P�,��yy�ٳ�ٙ�۴/��v2!���)(�n�F �}�˭Ǔ�9���|��s{U���C'������:�����D���gxz�q5��B�֏V��m�ϯ��4̳L���*hx�X�=���� ���D���|b�s7;��7V Z�PV�I��p�9��I.h��]��,�:�].��BuA�:�.�&M���z�SA�]�Efq�u]g��<1�Dg9�v��Ok�nf�gdɎkd�a�+��[z�m����;c�er�o{=E��&�Έ����E�r�����l�;E�M����+��(��8�x�}vx�pmnݨիl-<�n�6�ynQ�{F�!ϫ�}k����w�v��A��m㞎��H�m��v-{c���8��{}��s�hy}�~�V}|�{���A�N�\R�;�\�!��2��u�f"`���������a�Sѐ(���#��X*��\���v��Oo
�5m?߽�ͫ�}T����n|�'̤�o��]3i�m��w��ͳL�+�ݽ��R	$>e��b{���Maj=�甛l H%�U�Jf�L��x�O�	m���J&i�}���3I�k�r�N�I
�\5f�����
Q�ِ�i�5�R{��76�fҙ����٧���2ӹ���6��2����F��i8�f��8P�
J6�H%]|j�o�@ $��k���m5Oo�M3l�s>�Ž���-=�ߛ�2���{��z6��̨dp��1�i�#MB8�v#ZJI���O���I�e9��Il�3[��+B0��������	M��vųV�x87�ې��{1u����+��wGa�� *�J��"q��� c�\5��L�����m&ٔ�*��2�&Y�w�sg�	>f��Zc�z��%�L�W�����SbH�i�kMB9���b���z�[ܷ_K����z�dL�]��ʶ���ץN�j�W��>\]�.�K��Z/LI�7>�FYr�8�oo�V/���Ŋ��u0��@��@ƈ��"^$%2�,��X*i���-1q��>M3l�w>גͳĈ�|�o�/>���rD��H��T5�CK�ۭ5��#�����c�D�m�ϵ��fY�Rs����XD5���- �P���2�_2���A�K�u��>M3l�w>ו�l��N��si6��0	Lϼ{w8k�P�w����T���ZD5�S>��(�2�2�I�L�8nfm�fҙ��0T�)4�J�~yvͦ��S;({=�rD�D'e(���n�bD���z{u�Gj�`-=rîF�s7�l�~{��������3�ēpc�Vk��G�{�u�kiLǼ{vm�m�����=$��[ZE�}��0�#��԰D�,�&	�6�fҙ��Ʀ��HZm������6�f�L�}�f�l�);��[�Od��[/�qx|U9k.2f��8$��XF��u�!5�CXj��0�+&W��&��z�:	��a�]H0�*ئ�e�w;\��\nt�o��Y]��K��%;�ǰv��u;<�o�;js]`3<���1GIʋG�*�$Qɲ�F��wur.\ᔙTPT���@�)5�T린�}p�`�E�d}����II�L��e���}�0 w>�ųl��N���si6�f;Ӻ�Zi<H���ހi�D>����D#h������B���R����S��>ռh��e%g��*�i�m)g�ضm��@�x =^���#��!��M��Gb�4-l�b�����^N�ޗ���L5~w������-�p�|D |D5�=,i�l��{���Ze���fQ�W8�ԫ"L��ު}��d$-�i6̦s��p�# �a�;���l�M�)�U��e�L���N��x�A�|hOx��E����P�%�XD"�ϻ~h�M3)��ܢe;$�b4���C�Zj��]�U٬#�i�up1Шk#MVqX�f�m�$��^l�f�,�y���Zm�1ۥ����5îD�G�����Z�T�͐��H�yD�ص:f�Q;�;�n.����j�c����렬�- ��{�s}�і��H�U��L7�s�������A'�<湘C��W{h�M3)����J\R�JTFF���a��C�+B0�= $	u��l�4ϙL�}�f�l�x����ơ�"�P�ҽ"$4�N�l)պ9y�Yl;�'m<�\j�4�ᣝ�\�ߞ�����1���[���U�3�~��B��!�й�X��u(�e&I�[6�g�O�e&�I���#�D��B\D"n,�_��5���;�	�|�N�����L�S+<��UͳI�Rs=�,�W�`$�kMY�t����'
&Sa�li�kMD�iԩ�S4����ji��Dm����L�6Ͳ�������3�ZW<�|��9"JG�n��5�P�(UY����Uϙ��);��a�Jf�L�5mfY��@�Zs��ͳi��{��H��*�P�i�F��Ow�CZF��P�a��}>�|�'}Z�sl�m)���С��#�Y�s\CɟL��{�#���L�~G�cAl�S��z���V�םy��k5��7nL�)#o����997i�d����������G�.��,�	&�ec`�_=���PV�y�Mѳ�^��v��/d&F4	�&���x�&Q�q�n;U����n8nՍ�ۋ�rG�I�L�SN�Ǝ�ڕ<�n���݇��ܰa�eӥ�.�d�_O
���n������y���ٻg���Y����W�;t���8I��]��W=a+J��c��p7%�e�P������U&S*��g��� �0L.1�X�2�"&Z4ݷ���ߙ~�C��[��2v�m���f�FW�G���3`�]i�u��{���}�S���1�5xg�L���~W�4i��2��L�3L�S>��(���C�i>f�]�)!�c�z����L)R��8�sRͤ�2��_� L�S;�w�.m��g��߫�RL�|��i��5UCMB8=���D�l�$�V*�e��;SL��<�1t�&���Jg{�},��ٔ���2��,�{�Yҩ�L8\RHU� Y|(�(uߌ�6�5֍0�Np��Z�'P@
�f��cHF�+�"EG4d����i�P�=��6�he�I	�^��2�;Jgs��ş!i��y�,�h2E��=l:M�H8S���4sog��Qr���K���ݗ�:4�绻����}�ԑ�(�l|h|@dw��в��od�4�`���3g�	$i����ڱ���d&|�J3棅F����G���5μY�eo�-8j�;g�?������o�p���ώmV���r�hBs���tNe,���rʖ�{`�캻;1�����UⲓJ E����M�cwFI)�(�Gw�("��&X^/�KJI�k�ƍ$�2�|\�: �@4�9i���8��"% U�ư�4����0�f���r;$d!�I�V��2�&q�w�3s]>���!��R�P�-�z��@)�w^h�M3)�2Ke�Y���e&����	3~��tϓI2��{�*0�Z��i����b��&_��J�}�Y��m>a�W����ky}0a�L�P�h}~�cD��.���e뮧�vúq���=s[.v���CZ��k9#�1�B^����b*�(�IJ��ī�o<�;�4�`��.���L�9��Y�$���g̤�כ�f�,�=x}����\b0ۊ�H�4�❈՟P �HZJf���i&�)�3e�]�J�W����#Mc�x}��l���p�b�}�{jƐ5��NE��}�t��9�]ŗ9��?4+�Mޫ�ݨ%��.*㬫`Z��S��uT�WNspm�#����h͹<21*�Y�{1��S�t/6��T�90pA�#R4''u���3���C)�AAT�}L��s����9j�{��Up�]6$�w|(@
��ʙo~k���8�wuP��;�{��u�x��q� �����rc<�:��o��@
��7��Y������B�;���ɭ�k��dnۮ�y�y��Pp�i7:�B��郝y�q➷��{�}�c�^���R��?y��o��v�u��O� Ί -�����~�|^%8"��%��#N�gE�P8.�[ߚ�d���<���_}�y��P�"%�Q����~l���s/�G�ǽ��M��j�dvO5��P5A���hPb���D̴9wY|��w}O�x���|������#��k�|�79ܞ7ܢ]��2�{i�{tt��:*r�M�ZB��\\ɧ�W_/U[ܷM���S(ȩ��l�&q�(�(�"��H�;��r��rK9ь(�QEHC7���[e3iO��Y�Ƅ�7E��H^��,2jȆ��| �&o�b��ٶRc��4�f�ߎXk�P�Pߺ���02��F��6)�᫵Ϧ.�P�b燞ʑ-�{.�kP�v��(' h1��5�k�)��rͳ,�)9ҵ���L�S1�iJ=$ �4�e�9fVZS-�Ϭ�s!q��F�IEcH��_�<6�iܑ!&���}�ff���)1��stͦ��S9�^�g���%3�Rb�/����Q�7Zj�!���"V�i�Rc�2��3!L�b��Q�Y�"/�2�,�-7҃<2%"�sl�m�``�J����3��6�~N���Y�2ϙI�V���)�OH0�i��H����5��8��pD˂�m)�e3�%��l��m�W��f�L�S>�cEM2�L��o���0E�`�>����+�j�f�m]��)�����v4��t���R2�֭��c�O~(��Oaɵ�D>>�ּƷe�@��a�j�E�N�<������T��<���}���
��:\1�gTS�Z�9�Q�g�5)�QQz0nT��8[�q9�V�n����S�MTs�P�X^�I;VU�H�
`UTS��l�f�w�`J�j*�X �ѱW��|�?=�z�۟�[d��t8�Yxk{�9N�S���=��q\cb-�����bh��i�³�^����2	���z�yߌ1�^k�Y�-�)w��g����ݼ<:Η����}�ۈ�T��/w�ٹ9����W:�q3�ӓΜ�v��0jf)����8Wz�2VI�3N�h"�f�sNT���6?p�OV)�z^l�j�L�ݞgG�Z���	g8i�\�q@���n�e�둔}���y_�:�Z�MS��޶xCǵ�})����է|o�8��mlKnw6������6Lx��q���c+ϖ�#�	D����.��"J��1;C`�ٚXV�^�D� >j5�� �6M�6�޸�lS�)���N"�2Muj�-�$���E��hGv�egwJ�9�!(��g��>����NM�{�L#����x��y}8V]�����ڑOocN�D��kj|&�0�orX������+���B�p|����Ϭ^��^�w�
��3]�M��ݪ�U�6l-��{���P�+��� QiԮY�;*��1�4����=�H������ٺ��\8P�X	��=�	ܸ��Ggv')�?A�~;?�u]�b��:.'r��k��ts�W�燹�dy6��I��q��(��T��B:��`#�=�⇡�Ǹ痎t�p&i�W8;sɛGa�n����ۯFsۉ*���ݦ��\�zbw�:>}�\9���z-&B����M��6ӎ����k����xPw�nyr�x����M���y.Z93����5�׶��^����{�3���n�.f7���IT��Է]=*P�nOH5c�^���Lcn�<=�v{6�n�������S'��=���9׻[�qi��]
t���Tmۛ}̍�����6�r��	�؄�#!��2bkN�m�\@������K��/�����Z��� #��u���p���>�ܽ��|Rwo�덛Aj��[h��\<3�n9x��u�(�"�"�f絑8�[6����=��k�KI�ӜN˓�v��L�
荐��G�{�H�'�z��c��t���%��\��
5��v��E۷#�7A���ծ���T���h4�k�n�9G��
�<<u�:������nHәLm�rk�gGh���k�F��x�9��X�E�mv�������l��,d�`�g��n���h�P.�]�D�tw��	��qn�S&��'��W���`Q�u�p�s�]����{79�n�I��kN�v�8�\m�t�5�����>')�R�t�]��n��Cv�VǑr׮0����,&7�E�t�=����[��ݱ�4Xr�p�8�m�`�t]�3J�=�|y�v�������p�����v��bӒ�*�71�s[Xގ�z��s���v:��G.���t]����2���<�u�.��d���q���ۮRN|\c���닝�`�9����:2��H�/T:x��s���>z�=��i�g���Ƽ�n�Ϋvw�7`����<������nnz���Q�ۧy�4NS;s�:������[��6f1;�6��/^�r  �c�[6v+��-{p}��������>�*�N��'���sڦi6�z=d��7U�|��9�L���m�8��-���y7WSb��nI���F�\��i��Խxx���Yd�C���7��u���7��5���nb.��WY�Ll�f�ہ
�?ii%�f�=�����Y�tr�t!����Ǣa�4o wB�6I9����	���Rhz��w~���r�K=�qR8ӧn�P�>�<[fݷw���h幯�lӺp3�jV��3N6�}�(ŐZ�،ba���-�&gq"cÏ=��^�50��J���6�����uб�|Z�m��e�ы�y�Z]���x
ݒ�:���Ҧw��n�{0���k��V%2�i��Nl=�<[�d�&?
�z���;N�}�f��r���x�_'��L3N�\$��T��3 (�֍����/7�w����p��|9GQ�/^�O�^��[�\+�y���2�k��ٯ�7M_֬]�bA��h�:�����A��}G��FY)��eh�I�a,z��� �JS��3U\g����0cx�Z|=*���<;���������g��\�xQ�V:4ۇ%����^��Xl��F�����{Ӈ��e�u>�KY>
� 3�X��K��2K� �����\��';N�:�X��nL��:����FXJ��7��҆����=��ǎ#+:b���N9��!x��a"F)��m �AF<��De{nۘd�����(�%��,�\m̓c��ϱ�$׮��"ǷKi��v�uH���<�t���������>v#��F㑛\`���m��~׮�6�66�y���ܝ�=n� �1�y�V��u��gp���^̑�m���7<��6]��wBN��k�3�i�m�+�/د`M���{"ef���.�ؤ�;��۽��n�nJ$���W.lTX�m��G+��0�g�|�,ƻgF�^��ݼ�tm��'Kpn��d�\+`��vX]���{���~筎�I��ԕc�0׍Y���n��5�CK�ҕ4�M2�sE)�Bi�m�iN,�5f�
|B�2�I)Q�usl�m)�Ս���0�O���7߳tͦ��S��zM�e�e';Z�si�Q�Uf�"�w=h�:�a�D"D��i6�Lw�)f�٦S1\r[)�	$�-1�S3L�ZS7��EM2�MB��Q��'Q�p֑���![;�}���e�e'}Z�sl�m)��;�%ͳI���!!i��e,�[Xj����H�I��!���֚������e�=��u�6T�-6�Lz���3i���a�w��ig��6�G��I�4� �ceT���a�ņ:�;s�93�3uu�ܦvl��ۚ��{������)9FE�Cu�k�!���QZk�P��襚Kf�L�ד�S0$@!�e�hj�]J�P�f�9��*�(a�{��B'��4��>��>�z�|�¦>��W��H*i�)� MvHѯ�L�#�z�VKʋ�eHS��ӡ�Qu��MWdJ��24U���'�v"@�����>�&�u��I�f�F6,kr�e�����Y�e�e';Z�sl�m)��;�%ͳ���̴罋��@���G�ZE��P��,�#�L����f٤�$�il�+*m��j�}�kH�Zj�u��P��-g�b��ͳ,��$N����̦m)��}�%ͳI�Rc��K4��'ޒ �0Ԙ�P՚�h�_ȁQA��L�̹�S6��r���!I�S�# C7޽͇ɦ|��{��,�3�$�x�ihT4������EQPI��X$f�a�\�:7;]nn�Og�͵�S�mn7�{��+2� ���m)>"�4�^�"��l�R�̖�KB�Y٩GHKCil�+(��e&��;��	A8A��1���5w��"ƟP�	g��{����e3iL�}ݩg����������M��i�e���:�0�m�����5��ʕ����C�\�/X����\sB��r˸$>�?q�#�H�i�승v�8�8�ɪ7wʧv��܃�h��H�Vod8�s8��o��;�ˊ��*����%U����o�Bh
$���}y�,��%�D��9b�݉���Q�ڪ&���3i�m���۔m�f�I���	[��n]i�k}@*�U�}��R���m����YiL�S1[r[)������ ���fm�e�z�\z�"FJ$(��0�d?|y!�5��U *@�;�G��>e'�^�ͥ!��c���X����^���I�a�b.��ԧ���v�[��3^��띳ӹ&۝3��?:����p���	�I�VƇ�2}�%���;>*i)0����;$`I&���-1]���m4ͥ!\��SR�FLM�X�XF�!���i��!C��c���Y�4�e&=s!iL��1[��g!��2�g�äFXA#)A#FU��B�u��HZi����5[Ɠ���>e����ƴ�Cݞۭ5i��؏S�	��D�+J\�4� 0�I��ef�[2�g�8�S-�On���e3I����dHD����2.5�Q��3�694���s�A��p�%B�בS�Vӛ�h�ܚ��˞��Uա`�9s��~+&�H�s^\�tT�������Ŋ��CF3����E��UC৔�5FA���F�2&3CY�����6�gܮ�Y�S6�|H� =�ߛ�2��S1�{j\�4�e&;fVZS-�� }������M`ܣ2���^��q�۞{�pWfb
��tYM�v��i�
(���H����"V>5f�e'�N�M2���|]}��e&�I���.�ĉ�m�2��׷,�)6�;�O���a�ገ�7ZD i��{�,�x��6�2���ZS-)����Q�Zi����J�NI@�l�5����a1��8uV4�#MB{��oz��)�r��f�O��$��������B����3sX�}ޫ�"$))�*U�iL߉1 �=ם��̺��3IL�t�[2���Zf��b����5�Okl�X�#.��cMFm���k�Ͳ����FI!�{�*|ϓ�Rc�ee�2�L���4�f�h��1�ոf��VS>v�z�3
���ϧ�咥�t��ø��P�Uצ\u�˴'����T��Kb�a��5�^u�*g���a�[�_�xݗ#��ai$��W!�r�9cv:�\���&�����%{�6�XS�V� t�G[F�nlێ���Wk�磓n+�Lȯ�3��Y5��5A��Y�n��t㇫����K�*�\��Z�q�q����= [�m�Vw[�V@���%u]n5Ó�ϳ���
��I�կ�n.�G�nݸ��ˎ�{�|��6Jݮ���U�9��G��u�.�;n] ~}E��b��i5���,b�� �D�`��%�6J5�J""�ŷ�uY(�)TVk5����j�]�қq�h�-�ۏc��ٻ/K=�[�����ۇvY�.�WXj����ٔ�Rb���f��L�S?�nY�$` �Ց�#�%a�w�`O�3n����K6�M���+-�L��!l�2�s\�L�i�y��Ke0ˢ����'�Jq�J	�JjE���{���C�3��fSD����fl����5dCVj��_<T�(k9ÌSf�L��D���6�f���M�3)�Rb�ǗL�i�NΤ1 0׽��X��5��Ou����U����)�Jg/���i4�}8�I�h��%3L�b�r[)��Nn�J�6՚�,�Ы��<�h6"�Q�" ��ݮ�E!nE:ݤ����-k7l�6(�v}��w���Xd[��E�"���#�P�=���i�e3���Y�S6�O�N������-�Kg��3L�i����|��UpDm�&���5)�ŕfw׳3�MFBٸJ��ڹK㗔\�v�ϝ��ףq�z��g&z�L���/c^�yhELFa��\�����C�UNj)���O���-η�t��0�dX,�VF2PdѬs��ɍ�4kr�mQ����&�BQ��5d�H��#X=	!�e���xJ�e3iI��x��e4�LW���N�@ l�Ƭ��������.9V4�t�sڼb��L�S7����f���i�tef�,�S1_9-��e&+N"B�	�H�"�MC[*�P�=���0�`��}�&�e}��Y�g�0�II�kX�n��,�}xfP%�SP#�cHF��q�0,�n/h h
���<����̙9�a�F�r������`��"#����q�����3un����9�헮�Z�����}���w]���Q�d!8lˆ�#��v{f��|�N{m�76�fғ��'I��m�M��3fVZe��f7�J�u$@���͍5i��1 �	$$�i)��.��f}׷L�i&Y���6�E�l�	'̴����Wa�S2TE�u�P֑w؈u���B� z� ޶���>'�z��a�
�OV�;���XM>��]v�U\[��{�-5=#k+q򊵲Tm�0��<�n3�3�W�f��+����<�C{���	�U3m���@X�X0ʍL�6H�HB,����Z2b��F7+�E� �В�3��L�R{���5�C^�s&� �%���ͳ)����y��|�f�L�kۖm�Ͳ������e3o�	��J�ZF�}���"$'(�2U��L�R͙-�KB�I@���*m)�3���F��i���s�͆�Mi��+�$j^�¨�L�$l�.(M{uv�&u��t܋[�����N���x�^����p�|�,F�(�RRU��B> B;�+�"!��}�a2i&�I�y�S�Hm,֛>v-]���s)�bP��"�iHm)���4�� ��-1}�q�����=���e&Ф�u}�ͧ���@Y���^��i㐰�Isl��);�h��Jf�L�l�l��"@4�O���*m��%3���SL�i�D��_��\��5"�kH�[��B����G���e'}��,�[���&��{���%9�c-C�υ����e��!��d�v�vdnq��!\����F��F8S�����Q��ѫn�)Ѿ�TLvk�y���%+��Fs�sK��� i4Z+,Z��sQ%TS��ň���H#EF�d�6���b�lQb�أAX��$ü�E,�S4�-��q�FВ$BB�ƙ�5�f"%a�k�p�ā�t�*m�M����L�i�|�g��3l�|�`�������+"��4d�м�Q�77V�κ���s��Ș��e��=[�m���;�83梁�!G��7�>Jg;��*m�M����Y��i��;�B F��_i#rd#���#�B-�n�b��vkO�T4�Ƭ׻�fٶRwڿb��L�S>�w���z��_���.��'A �vl�v.�5f���Fd�   ��xEz��P��ޫ������y�fn"bh���٦m��-;��ع�I���}��o{8�cg�*�'p+�~�Gä8A#2��vo�Wm����( �����~�ݙ�z�Nb��4Z��� �w��ճ�"'/�L]�Ъ5��ʌ�t�9�Be�]�
�m��a���$o@�޺� �P�Ω��{4\cI���̾�L��g!oi�E����22�e��M�N�x���Y ݏu��㉊�.��9�n�n�u��K��B=�va�v�8���\���)�o;��7��qN��q{��;��½q^ѝ۞�����w��yؐ�A�u�.t�m��=�����bH������|�O��mN��c�/i��L��i�B[:�]c\�vql��x[�����\���v����PTm	��#X�Q�0kE�Ib�Z2Tj�ƧΪ�65v��F5X���}|���2�8���ݫ��QRu� �g���Wn��iؘ�]Y���w�����l��v28�"��:�cL���ٻ|\��(e
�{}��B�ˈ5��`�M�qm�l��v��4�����<�f��ڈ�ݜ]��<:L__/��Dh4�n�N�]��Ț�ޏG�}�4��_w����>�]��#"���qn�� }��t�Qbդ��Y��z"}�[��V�}�L1��a�KQ2�f���n�k��z��w�ͼ]��0�-��������to�;�\�v���n��^���<1��޸�.��������u;�g���.~~��`���i���7i�~�v����舿z0VP���w6Oz{[,����p�������̞*��/!|s����c���{5�{���:������y��{('&���詫�P�oM������+� N� �&n��U���ttz$zG��<X���v�@b���2�-�[����$��E�iAE"�R)�5��ֵ�糪�y'_0ghVP�_<w�E�Ɉ8Z�$�^����2s�7s�@AC�~}���݋��ۭ5i�C����!a4UcͰ��!I�^�Xa�̳��i��0�\�l��0)��7���i���}HDIr�E�-��B�a�io8Q�[4�B��ww6�a�w��`��4���f�������=HH"'vN�kc!�f<p�t����ͽ��Խ���_�j�ZYpN6�p�8j�Ogڕ4�f����h���i�Zc��⶟H&��-��u(�-�e&
�pa�d�HLfIu���"�0�	Z}B�������L�L�}��G7�l�-9�jT�n6��}}s�w5I��!b��L��u@0�5�x���T��}��o�	
��"�a��Ɍ۹=����H����9��ޠ ��^ox�~��M�'pnt���/d��NA8wh��_g��~���Af���C<\\����}/+������{�7��仧����wK�R6��g뽕�lA��O:��҅Tly�G������B[�~\�^�q��j�疣�`�����|1׎�|m�00.v�l�Ö��x�/so�[�A�Npf�OC��1|�]y)�%��8�,�S��G����y�$ŋۍ�6����#rΧ&���􁰇�V�M�jb�t�0ݨYy�m�q���|�";�ǐ?N��&Ⱥg�r�Z�v�T�<�	����x���h:���7��o�'�_�6�6�p�{e��wث+M8�xi`������(�Vf7t���N��]�iд9�e�sK��N�8W��87a�Ǧ�ɛ`���C�x���}0?p��:����T�W���sI;��O���&S"����92s�4����'|�g����>X�/R1�`���Z~�>7}����<��w+H��,���[�ss���,�Fwb��n�}�t�ӟ��6ژub�N��#7}�y��^��g*\D���i�*�'����Z��ť*��H}�d���/^3�禍ݻKvTP�)5j�w\�f�X��c2����Sݵ�n�b@I2Uv�gXF�Vdt*4hKu]���	F
��k��3�-L�_����'�$���yLǀT�����#��A�/��t*C�T/k��kCěT:޿,�����l�w�A��)��Ny����|����9ͧ��;�đ���������a���w�|Uy�C<�����| ���-����$'4�"͉s������2k��>>$�sID�t4�H�#5hj�xHAjk����S�����fg�@����x�HFۇ����剈��78��ë�B_b�� R|��ch��n\��:Svn\����\�S�7XA&B�Y+���X�ވ��X�9�7�;�y=^",;qk�wbv�f�K�Oe���l�Oq�#&���õwȥt�KG�nv���!Gc�9Ü��icIQ�n�dK9�o*W��L����X�x@�s�]VE��J%z?��)?<�0B#:7�/�]�%�����7p3/���G9����z6^���������I#�X8�z*�0�������5Պ�ck�S����"�-�&�*��:^H6�qr�^ۊ�v�9�>�3.G��0��y�En�	x�,���ST/Y�pck(�7������. ���{����>��O1Q�+H��ph�>!|���+�t�i'�nZ�S������Ɠ���������w����)�r,�k"�3�q�۾�O��L�^9���!�NΐX+k��2 �޷�t�z,�Ց�PDޜ���wS�^p.��f1B���b�u	��z z ��Z ��&˻�*1�Q��+���F�Lm�,m�Z6�Tk�rl[�h�y��mL!I�WusiHm)�t�R����)9�{���\�L�Hf��(*%��u捲�HRs<ԩ��4��g�EM0�t�JL���m��L�9��TY� ی�ّAcMY�49�ܺ�P�˯b�%O����M�����Q�Y�4�
�����d��"�`�3$ۚ���ݜkjl�՞��{qb;J�=[��c����w�Q�i��	*Bԕu�h3^�F	X�L�c��+L-�fY���M�L�C��n��4���|����m�	���K�f�l��t]a�|H��Ͳ��9�����Y�#���	Xk������c���~�0�!�
M]��0֚��;�F�l�)>��.m���|����ҧ��m���7Xf�,�)��ϰg��a2h4̆ƚ�Z{T #���6�������F���)1﹍�m����������?n�}�N�s�=��U��oj���\e�8j���췑u�9\nxWSQ�0�<��FM֤����v�j�:��rY�2�_�{�"F�`�3Qk���1lh��ljѹ�s�QFD`�0�zB���R�2�HQ���R�(T(����H�"�nQ�6�e>'�0ۧM�,�)�e��i��2����D�-2�Bp������p�x6��]�L��M��	"��\ᶝ�c@�S��alߞ�F>�H�l���|�O�>�Zf�I2���J4�f�I��b�L���g�l�OnT�6�O���c�B!NBF�v�|C5����~h��FM3l��y�SL�i�v�l��I�Rc��+l�x"��-��{�H�n6\ �V4՚�P���R��5��}��6����������,�!��Lha����)'#0��ˆP�HLL�o���
M�����m4�~KC��e���FKO��ZD a��:�Q8���.�a&�O,�b�IL2�$��|�Z6�he9�\�e�i)��p��>e�̴2������`�,���uֱ��!YP�xfo1xƠ�F��Brn.Vm����q�倊�g�ݜsen_9�X�95����@S~!&H���A�Yų��\��S�{�Q�n�δ�����1���٩�)�3��xҽ��6�v�ݶ�.�:�۱���n.%�i�g�-�'a^5e}�q�qF�]dmz�\pۃ t�DdN�)d���.ʝ/a#y�tn�o�˳s�v�s�n�p��9㇞}�GLe#ƭ�^3�c����ݶ=�X(Q��Ir�Τ�;�'g�Ƈ�H܈�����ﺮj(��Eb�cQ�*܍����E�BnW6#b���\�/}>�kݤ>+6�6&;*��N��f�AgO[���R\Y�n����o�l_k�o'��nٴ�6�f=�J4�f�I�7Ʀ�L�W�~�?|ϓ�Zv��e�Jf�G�Ի�M(�P���՚�P�>eJ��Aٴ�w�����I�Rc�}[f�L�)����i�$f��Z`�����АQ�u���"]�Ս5�i�N]=h�}�)s�ѻ�C��ʖ�����٤�-4T���"��P"�g�}�%�I�1��Q�Zi&�W�����o�����fS�/��tf�9����0�4̳�e�Hz �g��4�a�{����m�Lx�kL-�i��Euw�4ρ1���#��`K��`��M�6�'�t��&����jC��wֵ
8�-��>5f�48�f���k��\��)����x����S1���q.x$""BԕcCA���/�^�^�C*���u��ޑ�������ZwE�Jt�_7P�=��ܽ�%�!�1��������o?��/"��4���9�΃}���Lx+�MX5���E%����ƃ/�m�b����Z���6�/���x��w��e�L6b�Դ��!�{z����i@KmWZhi�G\=Xa�[2�l�(��4�l9�jTѨk�9�s�6���m?P"���{��O Y/���Yl>1]j[)�Y�}�SL4��!IʳՆy)�e3Y�艨K�F��$64՚�P��wjƵ��r����->e&<wնm4Ͳ���R�2��RzH{Ϝc�?)u�n�K�Jw�p�������w�]Wmv�I�n��d������N�A����{��L�S?�l��m6�Nf�����;e�5֍Im�f�i��R��L�S+���c����2�5di�B��f���"g̶w=ܣL�i����4�f����Ʀ��|�2Ӟ=&S8�2��F�xfҙ�S1��Ѧ[4�O�LB��!,���߲��-|���q+I/�T���2�s�ھ��'�F@|�];�S�z���%�9���`�f��������y�5��� ��E�����*-�4$2d����d�F�rţW*�lQ�6**�,jX>&S,��}l��4�2�=��6F�P׻=�$�q7j0L�cMCZ�!��t�驶V�<�uԹ�^똳�ưS4�!l�u��٦Rsλ�"p6��CM�u���"�!��5d�)�����W��4ϙL�{�F�L�)6f���)�JgBz�l�3)��&)���n�&'��E�;)�k�v��!�	j,\ә
�Q8
ū�(�PFK���Ց�N��V��i��|_4�f�I�oᣤ6�f���S��6�M�����H	���r�n�֑���5�̨0�@Kf�i�u��S4�Ϲ^�%Ͳ�l��l�a�Oa�`�m����uEaQ�(��5f��#���5k���6�H	�)1�ޭ���e�g�ha�k� ��N2̀���gER+�ﾤ�̴�);�=Xf����|_U�驊�6f����I&����JvX��6��t�9ǽ�dZ�z
A�����ڝ%�t��n�5�i��7<�d���;��f9Y$�S��DYܷ1��;��M~;�Tast�P�AO��]�d#����L�
L�܌(.��M��;��6�f�O����e3l���SL�i)����K�e��I�+���_��IQ@�Ba��
ܸݍŻ[�0rru{m�Ϸ����㞸z�?����E��ZѮp�4�/�5f��#���SL�i)�������2���ZF�P��M�E��d4ґ��e3l���SO�!l�[>�o�K�e&�I����4��2����F���5�Վ%� �a��Zp�5m���7��fXe7ӽ��hz@~e3���P�-�O���M'f�ҹ�gw��*2�p�H�WƯ� ��`�����WWi�Cj��"���&���Ii��De -���}}�1fON�&t�͟q����bɒzt?h�5�7=k!��h�~�[���@��
�D��Qw�ngګ��mᵱ�\�(���Fzn쳾�� t��:�n�������_uB���?�q��wn�6##6��ϡ��h�uɌ{3�?��m���8z�U�H���u����;������6�] �h�@\H�ι�F��yNޞ���s�k��͗��a�ͮ|=�;pn7�9��o�G��gl\�'(c�AG����z�+��Ltv�W�.�J<�wmõv�j���	�Vݞz�\N�4/k��GTE�˻K<.�%�F	�!����~s�ݚ6���R`��64m�H���y[��H[��`.�ƾ�/��}�m���q�ӫ��n�<� xz{*�ڎć%�Ʀɺ�u����}��s��m�����x��P�s��*��I�Rc��+i�3��>e����Ff��#�8Odd�!��F��P֑}ɞ�]i�N���P��rd���F�l�)>͟54� !l�
�z��i��P�ʺ�P�d{�Oa�L�7_^
��CL�������Ͱ�]��u���doG{�2��H���ɭ�ߡ1
fz_��2ٔ�xr��L�W�⥲��aI�w�����,���e(�m��A�L��;��a)������̴��q^ie�3L�c��Ѧ[4�^����i\#�3YÚ8Չ�m�հ��흟e�v����z9h���6����,���(�`�!�&�tY�����2c����5�a�5}|� ���f�i�ֺ��)�Jg����8������[��5di�G��ka.��JϪ��vU)0����:˔��Ȋˇ��ŕ������uH���Xy���L��WY���6WXl-ME��:�U]�y�(�\&"L8dY����A�H20��x�$TE<E�fS[�Q�[4�M�ε4�f���k�qsl����0!�)��Zhi�k�օC�e7�s�L�H��=�qf��Mw��K��w�@�j#M$b��3���&Yl;��ۚL��W{WL�'�k�� i�:z�c�8R٪�&Y��y�`��[��d�u�m�ٖc�{��2ٔ�?54�f������B�oAA1)�Q2YtܔK�Cf݉κ��;I��ټ��C��Еv���}͇��9rȤ�]|j�G����#�P���B�3,�)>�k����i�M3��^E֚���杇*	F&p���z��@h÷Ń�2d�s�V���;ٳ|(:��]��߂�@�N2i5ջ;�9�����;����?]��ۊ��߫vrt�J�2�t:�������S�kun�Qy��kb��5-�z��e�!ՙ�:��yS��X}Q���bc�\o6�{�#BB{��Sc^r���!��]$��w�鳓$[g�2	ހ�AT�Z�N�S7ٶI�{�{�8�M��پ��L�i�e3��޶m�ͧ����~n�5i�<p{�"�I�.H��{�e'3}if���S�1+�}�>e�O�i���Sl�i)�6�M���({,%�q�M���8R`�`CV�w�c��{r Oc#b8)\�Ⴕ�an��� ���H��ƥ�_:k�Vk��>64�5��sկ76�fҙ����<@d��O�h�Ma����g�3"nF�H<�*�6�f�I˧�M= �f����qsl��)1��=tͦ��S>��f��¬ЧXk�3�f�I�$(���媪n|�fҙ�S�˛e�JNf���"�Ti�4��6�N[<9�$��Q��rD��%�7�*U�g��}�'=�|u�Gݙ�u���!fyu��^!�/GT]����W��r�5Y6��x��T%����n�nƿؓ5�8��[��uϸ]bS���]=ݗ�{��Wk�1[��������ؕ�V��t#A����b6�wB��'�٣�X8E��0��d$`EçfȾӓ2z��2�����m-ٰ�uwf��������)�RLC
�%�of�=[��g�k�lXv�Tc]��K�[���Ē����`$B�[�b������Ų�p�
V޻S�Փ2s�:l'!����gvl�s�V�R��g�<���垺6�f�Ov����Љ_e�=N0c+
�BJ��>���ӓ$S�Փ��6����L��v�ݛ<Wl�L
(�A1k^�婢�9�����y�����ݭ�� �3��̂��.�"Z�C1�8+m�Ͳ��\�SL�i)�A����>e'̤ǯج�Il�)�}�ܳm3Zj���Ҿ.o�K]�.�[�?���Ss���8ɀ��8c�^�AOp�b�rjń���7���}�7Ƿğl������ѿƫ��h��d�r��E�,B�Xg�[5�3S�b��N2�%��}�Vr���E-�����ɀD��Ƞj���J��<M.;�5}r�\7���\^��Fp��b��o�xW,��	3_����T�y��Lr۷`�T��z~��\�q�瞘Ě;������5zwI9�(�	=�[�jsG4�Ȝ�a�v�n�R{��g���ʖ�h�9�6@��	QS 욭���r?\�iX)Zw	�}��˸����Dvn=2�V"�uv��d�����\�P��6�38:��B���οۺ�{cڜ�H�����]D�h�yR���ʷ/��WY�]�^Uc.r�_�s&��b����F��)��k�ש��
7V�moW���1k�%���=G��gR�F�4e���τz^��]�Ε�7u�_j�ۜGa�jɬ�6o�^�ۘ-�����>�j�=矻a�J�C�0���.�e�*7��ٌ�Y 1ݗ�ďxXqLyZ���mO���&����:�{[��{�Х�+&�L6�=��vpVv{��C��t��4��nM�j��a��g�οr2E����V+S1�ū��#Zl[}�՞���_yd�����@�'����+��IOQj��yN�d��P{'`����%��`o���ս��F�[aA�IliKLa�Bj�(+1�Y��{v��v�(�0����d{��>���'�gb��ߧBn�*Q�3c��/]�	Wq#`ZkZ�����W7�Ʈp8J�"Q,�E!���v�n:����꽲��������.z$�^�a�um��лY��ϲv��Җ环'b�M��l�ǫG�,���z��źE��*��:�\O�%��tlVv�G$Ud9�-�5����ع��kö���a��Yݑ�l���w=�C��|�8s��ދ�.']wn����]�=kmt�Wkg@��O�8:�s��r�V�Y&�m���q8(Żv�kx�u�+��Q��:�lI����;�;Z��k�#zkx���'�Oq�r��g9殇���w�ݯkt�vֹj �I���k� ����ݭc��[�Wq����7lb��#^V�ݮ{.���n��ֻ���N����7b���3��	�Ӵ�����{w=�ض,��=90�ڲ��6�up[f0���OR�w+�nt�rH8sy;lq�:�08�6���8�4�沏ngͺZ�5��S;Y�����5��nW���י�i��X1	�����ܯ��Ͱ�ne{1�:^��z�ێMٶB{;����K��b��'m�/�z�wD���s�n�[���.�6�E�1G�bE�P��Ñ���s��Lv�{Q��b�lvc��{V�ۇ�p�)�H&&.��U�A]�^&�on�h��J����`;sc4<��Fr�6�$�����K��p���QMpN
����]D��u��<�%�6��C�k���hœ��P�v���
��vvx�vD�r���'\���vٚ9@����!��4��Ő]�v�uw "[\�=��/$u�fѝǞ�Qpq���7�g,�p.�Zݺٶ�Һ4y�h���sv.2٥�pr�63̩�d7�VW*�]�s0a�H��N�y�X�;W:��W���/�{[�E���b�����/k�=�Xu�s�=)]�9ݏ8-0�lv�d����[���3l<���r��+�m�p���yڝٞ.N;�V�q�˨6�q�1�\�l��yxH��xZ�/��ι��N��c��ֻ��t��x���8�7���@��N=��t�e���ߨ~¼w!m��ӆ�si8�g����ӗ��b-ċ�˦v�K}� O1#�9��=��j�8�޹����0BH�N����(a"i�j��ټI�B±&��$2�z�D��6��}�L�ȏy{�S�׺{��&e��5��w�I��5lۯl$^c��ll:(���{�ۅ�:�K��R~�o[*�ոZ��3x\�-����`�J(=��N����U9������u�U�Fn�c��Y6G�8*���S��Cū��el��ý�<]����v)���'���zbg�!�Ri�g��/���  �/a����p;4����O�ç�t�;#�$�t���� �]녯�J�`!�|�d��=L&щn�ؑg�2<�����{JHV��'n-�vŇ]��y��Y�{�^'��,��Y�O��U�d6������/��f22� ɝ�\�P���^�t����͓�����a��5��XGF/9��,~ �Ԟ��)]|��J��C��$����Ý1�1�Í��5Ns�L�����^i�{^-�رzxo\NV�=τ�.,�viÿ8gf��\���>L%���ɯԾ����#}<;oJY.S�c���;�6eFPx�E'Ƭ�_�Ӊ�����U�*Lw{��SOMD\�f�=��~y h�XC1;��ܑ�;�>�h���;Z���܏Rk�}�<OE�e��.&��Oc���;���Dn��sq<tyϏgQ�2y�r.�ً���ڡ�Gt�d�S�m���5]��&�7�xE�y�9\�n����{`3z�5��Q�O<2��!9;t�h3�v�;�xw�����z�s�<�a���s�Z���f��������f�yFBȶn��~]���@��@���1��"E���wӹx��Og��EZk���f{g�����ڱ���C�L0��~�g��8Ͳ��L�m)��N�\�-6�Nf���4�2���1G���i�e�.����L�S>f�X>��e����5�P��ꍚ}I2�d�6�3���,�2Ͳ�ޭy��S6��g�w.m��t�2����3��ҌēL�5�CZj��pa�5��\�	XD� 5�5��p���B4����B4�5�����*�r�E)+z2;�e�={�s�S6���v\�-6�Nf���%3I�l��ѶS4�LP�zu�	�����.m�ͥ'����픛e>�g��=tϓL����sz�6�O�Z�sl�m)�!�[�}Y��)e�u�匶��7n�\�<�lu�Y�tf��6�8+�����u��bȇ^kN��̴�������Jf��_�ѦRi��g�v&�ٴ�w��Y�Rm�B�����O�M\j;�#i��Vz����A�*.�l������@5�)�p��ѷ��d�D�Ee�Pʑu�����������񀺻4p��T���~���5]�kv`*����E�m͋�F�M���y�'9z�sl6�g;]Ƌ�&���y֦�j�i�`��"�7#I �	�4�m�'{�eM0�e���LY��>e�=�cٰ�4ͥ!�׶Y�Rm'����*�)��nCu�B��P����ş$�e�k�D�-2���4̴;T����ޫ�F9rH�)�Y2�fS�q��vϐ̂�{rͲ�e>����m2�r����������IB35
P@�d ˎ i6�g��n�@�'�P�e�ñ��uZ�og\j������L��fP>��ʖ��{��Y�M2���f���|ʅ��*%IUi��ϻ}ni� �IL�{�|Y�-6���۔JfҐ��Ѧp%�������0�.4�,��"�H�"3���śB�l��o��l6�M��ޯ�d|�K�/�$��V��Ю� �l���ଡ଼�'�.T�^_N�ٜ
�*��a��g�^f�����I�ʝ#�Ny���{�םy�`qQATUX��h(�sn\��$�`U=��v��f�I�)=ɝ7ZD i�E����%�mM��2����&Yi�7»�4�M!I�լ%M%!��A-����|�#MB'���b*#A1j;H�6��9]ܳl���1=�ߛ�%!�S;�{eͲ�l��{��i)�e3�Pb�:SD�g��A�����e8C��'�ٴu��-��kC?�������"%{vk6|�g��Zw��%M����w���Ͳ�l����O��|ϙl�kۖm�kMB���_�N2����MCZ��f��6סO�����i2�2�_�ѦS4�O��a*i8@Kf��|t�O���r5 7Zj���/U3i�m���g�ķ0<Ƀ��Wk|n�5i��=�.�՚�ޅ�[�Fӎ$RlY5����P��9A��L�rqXj�C�;�7Xj>ƞ���9���VV`;��mr�z�~{�;%�MT�w9�A�.έs�slV%u���\Е��c��2�S��7[pI�2Gӆ�o��3&<���%c ����+��S4��L��3�	m�CQ��t�fS�W{sl�m� {�U�6�a�����A�L��k��e�Ф�'��w�
{7/n܍�b���7���3r�\����sD�`B�z�UmF)1�֍��y�Vk����=�il��)��;�0�e}\Գ����gݩ��4ã�;i�RQ�R��I��4�u(4�$CiHp��*KC)�W0��)�a�g�[�gI�R}}\ws��~��R� ����L�{/�]k4�{ʚe'��}���Ͳ�e=�h�k4�&�xL�F\�2PH4���4�O�����L�S;�����)6�O_q�,�i�O %����,��kMB=s���PĉM����i�kIL���u��ٔ�)����K6�f�L�u�Q�S4�O��a*i��%32�_t��8jd���[��&m��p]t�@l&�WlI}p�!�-�EU׷���z�'H�v��*w��bzS�}�m,yv��b�>��4NO���b0�5U�>;��c���I���׮��=
ёK��')t���S���;v��m�Au<]b��x���.Ň���v��^{�-1�^�N���y�:�L�f�����/<R�U���=ٽd;��k��c����b�G:L9Z瞛X�Ŝv�=Y��gyXθ�n���{=q��»��2x��ΒwQ�z�+��N�b{���s��j�b�*�Z���h��C��x�=�B�\on��=�ou�i(d�J��$�H;�F2��;�}=�9ۙ�_V+v��V�4@�f���1�R��f��\CǊz�-��Xh�bc^��[�[�c��(�4��2�����6�f�I�ֺ��
5񿕚�}����xzl��F#կeC\�`��*��Zk�'ȉZe3IL�{{�sl��)1��(�4�$a�5f��;�1�p(�a%%X�PͲ�ޭy���6�Ϲ���f�ˉ1�-;��m0�`�-��)���[��l�
$J�+9@!�w����&�I�_�YCIl�R}\ܳl��:H6����ϒ��S=t�+	��qK���ٴ2�e'/��&Y�����5�&ٴ����*i)%3����5�P����ez@���n@�m��ٲ4k�����5��[/Zv\OXߝ}v�ș�"&f��C�B�u|�PĤ����k�ͥ3iL����6zIi�e��#�<�D5�Bo�� �R4Q"=B0D!kD/X�{�iqf}���ߍ�\�Yte�F�����ח8��6N=�X��v��m���tv2Ś�U2��,�K�-��Uy�F���m��w�w�q}w���2�`����!��;�����E����-)�ow�6m
M���w7Hm4ͥ!�Ww,�<H%��,��^l�����)�!��!H���cf�6�Sl���Pi)<H�-�l�i
Nr�����4�͙�� i�n(�FƐ!{B����w�4ͥ!�׷,�)6�'{Z�siL�zaξ٦ͳ,2��<g�Y���.8�D6�������cMaj
�9���ҙ��{���l��)1��st֑���5���>�(#�A�%0�.t��f8;n�);9H�G��/Z�.�[y�0��r�IB�r�EG*�ơ��B=�nm�ͥ3�=٦��;�b���	��Zl��{���Zj��]c�6�DJUN+5���Roי�{O�ϟ���Zc��tϾ��|�g{^ܳl�m>m=�ߛ����f�"�{<��8*"�*S��Mͳ)�Rw6z��%3L�n�s4m�N~q�o("�>K�f�ϖQ),Ƞ�L�zM�w\V���GBn0�Y��O2�*sX����Z�xTg!�r�13�w!��NC�%\�lV7��$D ���!0#1IhQTX���x�s�>��	���s��ݛ�K���o��
�f��)U��}�A��g���vlp�F�4��H_fZْ(9��)�@TLI�����$FbŞ�>��x��B����#i��wkwvxU_H��F7��[p���\�����7>����ׇyv,�n���m�D�,0p���c���dP�8�TuͫJr���#ѐ�"��"7&H���QlH����P87^��ΜY�z1�w|�������1bz;"�gޏ'\����QFX�-�"���ݜ�9Yk��eK�p�h|��/�@vA�%Ip##@�+ow�P�<�ݙ>���[<�uͫ�<����ϭ��� 2���*�QAm{�ߞ�`�Uy�؇���^y�0�����f6k���<��1+T~0czW���������EDFq1�&2M��.�R$	 �5>��ݜ��l�d�H���'�#0���蟫�-;i>m}5��Z������FD�0Oj�q�]��]\`K�Ƹ��b��� j���ny���kf�6�P�H�!���yߌ$d���gw��'9N��;KCio��{,�F��N��"�����ȣ�4�3iHs�ܣo�>���μ��RJg�{�%�C)�R{7Ԡ�z@�M�����d��FR����ƚ�4���M%!��o�7�͡���̴Ǵ��|F�S�����<���}!��p��[=B��;��J���i�G��#XJf�L�|si��'dӕ�ʛe3DCK�iu�O���e���L�5ǭ�e�oX��"s��Q�>g̤�o�f!o�[R�֑������ї��Z�h���u5��n*Y��E=�;�wr��y����p��pŎ�s|1���.zy)B����HR%���V�n�c���\�����2A1!q�*T$�wp�kp�kn�nv�����'��-�+a�=v8�mv�*�1���q�`����9v�$YgC�ػa�Ȧ$7��B)�P4����^9�8㷷fۋ��ڮ��$�ݮv�ٌ�v���]c�WE�J�t���&�'O9Jz�����n�u�<��kv�Nu�S��n^{N@�Q����7��k8���f+9�S�آ*�Aa>��F���y�3 ����L��ȡ����+�����kn{u�KۮWM��f2���G�_}�#���RSNѭ"�Pҟ(0՚�)>�ڕ4�����pޛ='��Zp��ϔ�Xt�����M�	�Vg)g��m
Of����Cil���ҍ���)=�h��S4��+�͚k�ƫ��W�:��m�fR��U.m)&Y�x�[6�l�c��KOI�i���s_u(�6Ͳ�پ�4�fr��28!@�*S�5*�Ma{$KOW�N�S4�f+�{�6�3l��y�������}���L�5S�!Лe�JL8��5�Y�5s�� �ZkYO�կ56�fҙ�]L�3I�R{<� �!�":s��RH�1Ue��2V�G҃�F�Z�v����n�xN��"H��(�, �q����w��f�I�o���Y��s�S��^ f���;������"��O�1��	�X�#�y������׿G�F�Ɋ.�Sbf�;[�t�L�r=�[��Uavr������whj���/�ڳ3�g*��{�_��;"g�� 5ݷ4I�6�[��29�e�K�8Q2�L��x��m�M�s��J�=CV1Vj�ҺP�F�*"⩬\��)�Wq��3,�9ԣl��D���κ��)�Jg��5*i��e&�={j��j&(Z��m)����2���͜f��R{��T�)�Jf�ͺ�ͳ)���g��=tϓL�)��)�Cjdh�4��P�����T�%>�O��ܩ�Zm���tR�%3L�b�=�ٶi6�'d:�W�;�e���-v*vt/n�<�s�t�S�a�n����n�\���^Ÿ��V)J�v3�����%3���b͡��)1��;�������#6�I�;�74��,��ˏ��r����c2ͤ�2��nT=$i�JC��ٶi�a��R�L2�}��b���>5���(��!	�j\4,�l�zz��l����sL�������������c��%�v"CU#K���f�E���En�)�zg�nY�#���/�����[�~uԧ=Q8������]u�a7}ɀC���W����o���G2�^�YW����ؗ��^:��C��͹V�A����l5���7���u�l���gbp'��æ���!�����܌�|��r�j��E�t��n� x��;��umtd8�]��Ggv��5%1t�x5�E\�d[Yf�������ʜ�O5�=�6��*�Y���`N+�R�g���z�h:a��继�轮����0�/V\���M>y�Y0J�գ)��D� gk^):��� v�'��b�w�� Rd=��0fu��,��Z����:���5f6�'��5�@ݻ�z�X�4f�(�×k�ʖ9%Lj�'A�*�G �ۡ	��
����%v�[ť>��r�Pt�,��S�S!��C�fq*�W�+�K �Vz{�� uu��ԝ�t�O���7l�WNx�k�z��i.i����<�|��pzf��8WcC��'c�\ح�*/�����}%�2/��}�ϵtܒ��	��5���휵~9*���0��͇׫I0�ȃ꓋{�5�3����zn]]M��{:��Oj9��8�C��]d��<����u_fz3�=)�>��7��	;��y�n���bќ�����?��X����'�*{y�A��K��ʨRqЂ�z+��H�Q�շҴ�����n��w@�Xؾ�*]���9�v(�so��m��c�ѥy[���ܥg��� ��F7~ f�,9�^{�x矖z������1�OlD{n���^�:��l�9+ܽ�g�yEz����N�,��W�(�W��+d�u�ˁ	�a�j�5���:�3�{�+����q5Xj��Qt��"r�"Y���3�=��9��������Q싫����ۀ;�W���ā�[��GU�3�^���r�Q����>����HFlL�Ċ8_3�+���j��^tǾ�a�Szj��g*ɋ�.a9yQ�"U����v�U�7���$aZ�Kl`�I�r��t��Ɍ!0�\����m�~��P?w��e�?4�� ���BJ<k<}�4Ky�V�c�������S&N8=�+�v�y#�/�c��A���kI�`������u���T�{��c\O�0��B�@zh��G;}=�T��e�)p��6曚P��W���NsT:��n�F��p�_�=���K�Dκ�|;^�Z�)`.=��G+���<!\Н��Ox�����\Q7��x�<n�.Q޷�N��p�֘�0�X�sYt}�Z��t�ql�t�Q�\�iՕ��x)"@kC��9M�4n&��t�1�p0s��/�A�.�|�B���[=�|=Vb#�$}�/����{Bd���BK����X~�����)��+p.�G�n����1C�&$��w3`cH �TFL�D�Bidc��d�-��	�=v���4�L�}�YK�ٖ}�7��K���,�,i�5�� @�aʓL�g�����m�Lz���0�i<F@
�}��֚��.���p���c5��sl�m)��5���Zi�� �wD&��kMCJpyA�����9��������%�؈Lq�LB6Ԏ�]�	�2��Y�m�3�6[��p���Z�q�qd�$m��Y_d|j�~^�kH�Zj��wm�f�I�{��x�4��;��H��F��G�4W\i�a�SL�ҙ��1\=�4�4��%��;�6�����wn�f��m����͆��u���g��J$�r��8Y���6�'3�y���6�ϳ�e(���-9�u(6��%!���Q�Zi
LW����D�r��Fe]i����,�}﷌Y��e&+��l6�fҐ��rY�E��߇8�[w�����x��Ź%���S�w�=���z�~:�yQ��.�	 ;V�8Wt����n�kVӷ�=�arS[1o������"���R'5�o�v����Ν�$Z��ň�j7+����T�&�lF��@����"�i�o�{���b��r�m��e'3}J�Jf�O�7ø�l�m���:�4�f���sz�.m��e'dj��U(�8��a��9(�n]s]���yˎ��ٖl�v
j�	ƭS��ې�R���x�|E����b�CVe&��|ٶ�Y�g�ԣ��٦�����i�L����m@XA��Іi�N}O
�{�Ͱ�{[�sL����;����7�U3Y��'�	1
*0�l�n�՚�!�?,�0Ց��;���Gh f�<�[���m�+J�fFeDJPA�8*����l��w�ߎL���ϫ+�y>���%�B
\:vl��|�fO
���̙=���vl��Yx�X��Y��q��!�}:��w���_NpJo�36���ːsTN6�Ӊ�5�sL����EfLvp-�~�۩�/����glZ�[�C���v����z79�9^��ԉ=�[IVu;��fN��c@r1����C�h+��7��E�n��0<�:�k��ڸ]�c��;�NW]$�4<���{v�9�$�T6z:���v�p��CokZ������1�tuvo9&4m�e�xKb�Nޒ{pt����0󌷎�[(q�&�����/N�W�uԒ��Mm�r�=qr-���1cY�L��
�&L�u �I�D�i�D &�;$m�%D
��N4�c��h�ݽZ8}���=]���y^��nm��b\,"������{>]YY���g=U[�w�>Y��=c�\Q�ԑ2��x~ӱٟDDS���+����E���oFw�g���G̨l��t�u�{;��"��N���?ee˝��ѻ6vy.�Q8�B2G#���������NvgN�����̼�39��>�6���$�rD���S��Z��z=�8�Ӄ��[���2x /����-��A�#d9[Fs/�^P�u&���狝����k��[�v�%,)�-c!c�s����_O3��$_Y��/s]����öWX@q8K6\bٰ���79�GX������Љ�u���B�\�{mCir�!.�����㌼���{o��Z�7��.���㫡O�h�Ǘ������;���62����鱊�F"�M�`�s�b�1Th� Q(�	�n�F>n�z���8���;B�7-w���\�Q���,�ḋn��@���>��M���{76I�gA�J$�r��H�׻�(+�|~ٳ��+2�}8p�g@�b�0�l̆x�>��L����2V���g�U���Ɠ�uZo�n��s��Do�JX�9W����U䧵@e���&fu�;�^;j�)c��F��bۖ�l���)�`|�5�������ٵv�+��Wu�v23�:|��J6�0��p'ow6O��� &��zu��/,������v�۵`w����`4��
��g��}˳#1K�_����1�$��ډ�������i�_A���\�=5��-mU��	��}Z�z��V:u�i,��f.�fP�]=��/{f�䱶�!����!�"Ma����/-�X�ѱjأI�ڿ*�-�)���|\�(���}��3_�v�'3'f�BD�jI��P|~[[���ә�"�ϖL��U���%Ⱦ+��p1P��0n͇�����=@ɞ#]��^t�͟#����;ѝ��XYj !�	!�)��,��ذlm�������v��:+g�:�������!0� ����5���Aת�/�C#j����g�����;�H��-�ap���kݜ�Ν�P_��}��y8�qd��� /w9��h+�Hʑ��u�6{�C#1b��,���5Zo�n�82��y/3��B��2�UJw��{����#"�U�#+{���r_NUY;od���l�A���{�n�d�X��Tb�Ԭhͱ�7t�ډ�u��|�&��W�����b���4�n3/p��� �E\�6��E�m��Q��&!��!F��EX�.��ۀ`()�Ay��^��ĻԢq��d& �G����HW~�z������U-�S=�lt �$a��ѧ^���8�L�%�:;i���\��ٳ�?���������L)-�#��Sm����?6~A}�s�+�yԺ�}L����n���]]�PY9��������#��ઇsF���0X(&��|=�d,�d��DER�w^,�:�UG���ar@�q�:wzH�=�K��C��2{��F�ފ�W���~͒x�G�)�*(���{���ӯvz��}��{8��.ե9]�����6��ͪ�B�H/�B
����ӡ���h�B٭ʪ��/jLL�v��1n��ݓs�W2���/]jc_Fw;B�dU>�F���u�q��.3��s����KI�v�u�NR��^�lzmm����˹�r���;8G�2�=i��ݺ�_N2��s��ќ�gOl�2M��ԗk��/q�gΦ�V�{!ȵ�s��tX8�����w=��s�޻��e���Çvnx�gc#pi#Z����]��m8�K̢�la@��]�հ=����%�=�c�7*�Ϝw�{����;��{��lb���Z�F�1F$�b")(�F
��mE���E��6L��������j-�c�������5&9�9ݶ ��N��7i�����
�ʷ�Ow�h�{�;��l��Α�i���0�'�����^!1)'�����{щK��Tu��v��`�]���4.�}>�"*6܄$�P(��M���_�����_{�쏟��NW�%	�� \m7i��P�����dWN.��͙;ލ���yN�h���L�U�{��>{����~"T��(Ԓٳ�{���_z=k�X�.>6�����w���~�~��C�r��ۇuW�:Ō>��]�u��x��b�tKvv(]ظ�Ka)98~��呗�t��e�_�m��1oY�X�P�%Ï��{�ڋ�U�9��s�ne<ז�*�v*Dwt�<̘���z�I�g}]zS��!ss[�,f=Q5{Q�)�m��Z�����VB,�0QUb�)�Qh�b1�QDI��PQ���ڸ�Ɗ(�W5҈h�}��[��߇�)�̇�U�'}	��܉"%'�ޯ_����� ���n����<ϡ�A\qƔ��E�vj��Ώ-�Y]ﰙ~�;�����W��v�}}-y�m8�M�(3��d�h������t��<���f�����.8pd&@�!��D��lpI�N���(�k�>��4�m�K����"��'�w�f��-�q�{���N�n���7� �b�Ɗa�5�9�b�EVO��v��/���x &����qC�SI���	���s��-����Q#��el=�tW�]z�h�pܜ<���9�J˹ 5�w;��E�Q2��)���nr��n�E���ݾ��?6�M[F�d�Z1(ZZ+-$X�Pl�`�ؓ~�wk�$� �j��?c��U�.��l��8Qb8h6�[�� D��l�o�������̽���lt�c�� z�.Hn"�:@��:�;��tQ��UXo�v�}�r���mF�98��Z��� �n/<7ll�;J�f��A�۫R�u��)z l�����,�{�Ù���g� ̑sÙ3��}���A�BP����>�Y���u�_q�[�/��
�;θ!,FSBF��$�9�y:|s\��K�W�����p��e|}�"%F��R�@�s%�@���a�л��}�q�3����ְ|����.;E��Jh�ˆ^r��V:{ ]��Z��0�R���.�3(�Z3��=[ea�Fxk3h��rq|�I]��\��c?`���w��YH�)`.�1�-��b�,�d�Ѣܫ�}�܈�o5#D�kA"�_O��xwޅ�M�p(a����UV������K7�w}�����2D�NB�����D:�t]_��_?F׎zH��e�Se�^x��0��$�:��~}7�3��@�2��Um���q��J�Rtc(F�%8��Es�~�Pм��1O�ߕ�߽Ń�w� �s���P�%å�k�ə��Њ������������� oBEJ����Þ��W�VE��X����}6]�����ٙ�}��NH�QF�I&�]�����?{����V�B�nn��ϗ��i�9ΛZu-���y��9V���˚����c#t��Bd��bX�;_��c�E�㟔��^���Z|�&�f�[�q3J5�����"�����k�T�Ńj�,�Lѐ���������s�^��N�ظ�9�j(A;D�R�9{���ܗy.mJ�ucVI�)�aP������T4��$�����}tX����[���cg��&ۛ���v���T�>�8E�j��\��~�WY��eS7�<�}��B��e�1/<�Djɡ�:egN�������Ք蟿d�%��_"gG$�A;��wx�C<J�G7�]��4q��J�g�KMB�o>��{!,#�K7�.�!��pm�k*�.�.�O�M]�?Y�n@7���	;Y_�7��o��5~�rɧ��C�܅������m�N�W��I���-�⟽�!):v��1�MK:�3zE���偹c:=�vr��
�3��������C���n�Ź�N\������)б:&���!݋���ApC�gn�]_�[�zg"`[�m5w��fc�7���j�-�a�H�V�wyh�l�N�P[��0�y�G��L��Q�p�Q/�n3��3��>�жe��5�.�X��u��/3\�������30>���G��̬�S��ƭ�Ba����nN/ۋ�&c*z��c�{�n�v�r���9��!�n���{��u�̃�cL�X2D���CcUӓz�,���|lG\W4M�Z`V�o���ԉ7������¶q��8��x6G����:U�?���t�6���� մ,,�s �2�Ti�w�
[�>�����(�P �0�Q���4l<�D��h�#X�S��s��;�����Ė�S���l��v܎q.�v����A�q���g�wOms�a��h6ŋ��P�����k����i�w[6�ӝ]vsv�!��c��m`�-��Ѫ���F`͙k��;Hɶ�ݽm5a�r �@�j�Gm�}!�sژ�p� �m�!jN�+p	#k�ݮm�[Wn�`�&=)�k[��2�6���mk���u�v�|.��s��w�a2pOk� E���z�n�u�v�nN�r�Ω^�8-���UշG:�qD�׋����;!Χ�E�'k	�mIã��#l�V���i�d.�suuD����Z0�xw
k�<'M��e��hݳq��V��n�6��; '$s�f���v�^|��=�A�eX�l�n��2;�+887�'���q���DϣE��Şkkjj���\��{k�P��>��}�W�2�f,���]n�z�'��s��u�Nw=)�o]�m��G�ٞ'��p�b����m�����ݬ&�F^/��<�e��k�]3�ni<�μ�A�Ӯ���Y�x�1�:�ӭ��.�ݝ����37nx�mz�Ӟ�v��mbw��+��\v��u�sln�C&���7]x�B�Ƴ�k��qC0����t��h:l�og�܁�6��{]�[��HlZn;{�Ee޷g�k8�ѯ �v����[Ws�Z7�Wm<)�����5%&ְ�k5^�EƵwKS���qOlݚ\�m�W��n67h6�ڭ�q3p�ǫ�1Gkwms���kix���L+�{K8K=t��+�)%ϰ����P��ݞ��z���C�:����x�[�x��ѣ�{s��<;�u�8����_/K��7�����Z���W�y�E���-�����'W�=β���z�X�K��0��\�޶��ɧ��77Gm���ێ�X|��p��3kG\b�#oH��]����[1� Fܫ��n�V4���v�v�)V���Gv�[c9n�]t���\O֣�oAPu����ՙ��%�� �!5�����<�;��#=��#��39n�%��i�ͣ�d|�Hq� �n��z`1t�x_L"c���n���l�p����P\�I��������X�� 1��ԥ�I��c����!g���צOjtd����f�R���cp6ՀD��,�VG����=�:�R>��ϊ:�;Z>�D�I��Ə�X.Ń��f[^շ$�g�=��J�܅��zOOoF��Ɏ��n����ڱ�}�뛏 ٜ��qc�<ob�rުx��n��Cl��.�����V�1m���OHp��-�ۅ��@���9\�Yg8���{^�㻻w���sCG""$S��I�����P��x9s!���IM�L�eb¢#�ub���qBC=29�����XN#15� ��a5����`�L@̥�����N��Xa�$ɵ}r��Yν��4�!�AEO��jb��r��T�3�6>�>L�l;���&�o��'����6ҧb�sW���R��������d���� ���jɫ�7y�����q���F�%.��'��PÄg[�F����i[wM$<�+;�\cB�))��yz��o�0�nQ��k0&s�ݱ8���D^�S�jl�-`D�v�yH����#�d�m"��ב=��D�����REXspst1�H�Cj���X�|Z������	�Z�Ť��X��Xٖ��6�Y��C/"�+=�o_�.��ǅ�YL��i�abnG���R�C!ҫ��S2��]��Ay���Lr��U7"��=O1�v׍՚���D�譹��`+����[Oel�!�C>Snږ�x���\��:9ɴlQ4��v=�8�>�"n�V7n���c�h;B��Qa[����݉�I���'6:�9�Z�i���q����U���T�Wn��GY9�M]�[�m����vݷFלJ,j4P��\��b-d����4Q�χ�����s�{����8�����&|���v�����\��DT�l��Qm�QTI�}�|O�˶��d���h�
��;��J�_w֏�(�F""L(E%x�K���nhwl��C%����c�x'd&Q2EI��ɗ�����問�
�y�y}�k��վr���T��i���ފs�`�ُ��9�|+��9�j"�v�]o�4p$�-�V<g����k� rǭb��o�[���V:rc��w����a0�F0[Omt���v6�kth��#;6y�ݴ�֘�f�z��# #"��	
$�L�_GM�/vȋ�~����6l<���s^��M�Zi6�����'1l��ͼ���֮.��8E���Q|'��VN�������qP������F7u�J�.ݹU\t|(�=�X��Lml�)��N��K�t͸��شF~�=���@X��%1(���`����P��D�A�9&#c�2�w��t�����P�lߏd��А��Q����z�
�X���̿�<��|����~��M�$AHK��� <}�ݘ���o���fp '{�е�=�����nQ�(��̼-G)���z3�86��Q�_p�L}���.{�&ŨLd�RFb�	�#�:�綋 �Ҡ��S�Q;[l���q$&H��	�`�ܽ��v�1��tM�#>�Ͻ�
�����x 
0�`�Sln�|D�O�}�����]l�,���Vp
ٷ��%v$�1�d��$�����f^���{.��r�$mr�-:+v�CQ�̵V�x���^&n�y�&m���B�(u����¤@����`g�5��%d��;�l�\�Ϭ��Uu_*�!���Eb���0����4��s��w����&�E3�1G�G��~��ĺmO���H�P���ݛꪊtyd��s9��˜v�E�{�^.��}�d5	�S&oy}9�� ����j��ݣ��}^�0u�J$��L8aPG sm����^�v]�mq.͇=�)@첝4n����a��R&�I&ݏݿx-�ew��VN8��^�s��2�=�Y
B�	%(D>m5Ҿ/�謠�:iQ�ۉx��啝�@����g�R0�bB"�^Q�z�FgDE�:��(ܽ���������m�"ɝ�{��Y6l��ve�u�u�B�[U�.؊����}�Sx2�Jl�־�Ot��p�%�1���Q�m��ꂚä��q���JU1<�ÃrYV���[I83���~v��*_�:��IҦA]�w�;��D�r�u���	 
H�RI ����
}c��>���~U!�F�qHvnϑ���=U_<��d^̙��q�N
���I�x�{nm��z^��7�7c[Z"�֊�62�깖��y�jZL��m7bݕ��7�g���1e�[�33�������ȯU*@�$�.3-�l�ٲ/fx
�|�Ўd���l�ٰ�w�7�U�]�=V=	4�fL3��8��;���n������m�>���x���T� �p#�����V�g�>��k�,t�g�����w���g���A	p��1�qX��{�v����ًw\H���[Bl�W���.7��ĉn.;����b�m�m����כ3"5E�A�R�m�Y6��Y�!��-Ӥ9]v��|����^�Z�:>dq���:EJ��+F�ݾ���U��gZ�Hm��]�y�m=�6;\���E�tc�u��u�/7R�b���
��hלv �pa���E�v]�d�yMۋb9e�Bg�6�Aٜ6�]��/�9s����[���7X�ӹӳ�,�*�g{��v��휚�p{u3���ȧDv2�jF�h�v�5���l���w+m�s<;���Z�=]�p#����w��{חF$������ ���u۾u�w;��ۻ�M������ն�s��0�qn�y�:�c��>M�\&H������]�y������� U�����Uu���|EG�jӝ�]�m�<�q��D�2c�9�� n�w;ec�y��n��{�Y`�6���ဨ`	TmF�{�l+Z��ꡞ=�d��s9��9\�@LmE$���+t�P��{��~��ݾO��3��s�����g�b@X�!%û5���/P�0#���唭��2������RX��z狛�#���f9�0^�9ͼM@j�ً��Ik.ڴ�1�,l������Ͼ�ƅzjr_����ݪSN:�ęE �J�����3�~\��imoa�����|i��U��w��N�'�a�;9,C��}p%��yX���΍6_#v{��_:-�s"k�����P�K�z`H�薻���e<�����L�i@)"�B*@�-#F�!&�������k�Dz�)�΂��d�J$�%$/Y���v�)ݳ�ױ9w��B���ޒ�ABĄ&$A��� %G/^����+�z#�^��2�{�rPH��� �(��obn��ޥ�6e���ٙ,���+p�&mW	�ɍ�K�A���-�N�+c���[7��7��)f����Fҍ5��?w��g����ٌ����_��[W����D��E7���}ٟ{��גGSٻ������б���b
&�	�>ٿE�fK|�0#�q���l��0c�n7&-{7�Sx��׷��vM�׮��f�QJٳ�%T7}����dS�3�[�����}�[�=�n3�>53C�(��"m@ |$B�f�g�be�wI��\�AdX�p���q��/�9��k�p��)��1(�u�����[���Õ����=T*.�2[����Q@�T�(�Gw_=}���c�燽����n���}ř���V������i>�ۣSm�6�1\v7k�\�g�=)�F�v�g����
l8�`��2��矆c�yʥE�/��F��WWP�6Gt}��� 1�p9�������P��黷���x��.�T�A߸�P��%�D�)O�½U8Ӂ[��Y����ꏅݜ\z�,4��	2mF�w�9�Y�׏����viU=�Ѓ�˴���?U�MP�	�T��AV�q�om�x��ר}BW��}7zyG}k��}i�Q�b�`\*y�*N�ɴ��s�RM�k�AN��+�PI`�d�ܹ�� � A��<��U�=�����-�#�����?tw2��@}�9���E{��+_
�s�/!%Ȕ Q�dK��\!sf������)ʼ��6ykr��<�S�ٷ�&A��/yH�t�]���P��~�O�^>�����ԑ(T�79x�>7�C2o9�S���Ɍ�q_E��oA�12La����}���,g���_�Ul��2���UE�tAy(IIy)!z�� N�xn�e���y9���� ��w�}���%Ȃ�B�D���o���߅�����V<~^��k�tq:>vn����TI�wjw�I��H���6���ԛ�y���|J�rI����T���P�U��%_�s����;+��d�ˡ�ϯ��cҚQ�d�����$����m��җgsc�����6���Ƭ�w1�#���u�n�m�x�o�nj��-�ϛ���z��[�1m>�g<��a웶�.��)�tU��'��\�=��b�u���y�� �6��j��ukVc���^���p�D�t�pl����t�XC��v���ڸ��[�#t��tû�2yq�w���{ϝ����Ѥ�� F"���ĹF64[�<��(ֽ���ޛ�~tm�ٯ4�ڝ�N; k�go`Jn&��Pչ�Zi�׍W����~����|���C��ןG�z'j�����`�� �(�N)���g��6����� �M*nz�""�b�O(�	 % Zn,�k�x�o9���[���;����Vb<�:Xu$(# �8�k��K�ps+3�|��:(��/}�k��3�"SfQ
ffd!u'���o�z+��ÆY��Ɍ���[� 	 }����1����.ݻ�A������Qgr:�Y.�9,�[k��h�MGQDIB"`��s�~���M�ϧ�/\8}��f'�_�3����)�a����:s:/�_�_��� T�|sf�g����}�8�ioz~˛L
�8��h?�����,;�ޜ%d]ӎQՕ�;�S�G{spN��̼�a�1��8��0�D�p�sWݫ��vm;��T�j�,��o��fg�{�ź=�����(�r�l8�O�5�x��c�w:w|(�Q�n?��9�C|��P��%�D�ɝ 	��kw{}���{�����<|s-�]�0Dр$�Q������,׀�{�wQ\N/�~��gA��[V����jk]v%�,ݰ�Z5��i��]�8�OPD"���WXh����ɞ����ކ��|f����;�Pd"%û���
�o�s�3=ދ���绻�U���"��
�7E�ky�{w{޵b�Xג��gmɡ�w�;��Te��&��]�	�\w��@�M��U�w��p\��^�pz��Qt(U��J}�k���y I%4�b]�&����'l����l:��͈�(���Ź�*L���Ծ�;Q�}�(�����������a$mӔ=�j^Y8O�zt���QnF��<R�b�=ä����˾�7�j�a��:���w�w6�R���a��eD�(�'���`�L�N�(�����d�����w�y�	�&��؝��Na+%AQ�ri�Q�Gg�� n���~8��x����BT?)�t��aY����>"�����za��`�tn���޻�^n�z-�vn�f�|�ƻ��[�lw@�7�D�W#���2��[.�\��78Gs=NT�c�"��3��Q�Ӵ�dH�:��,�ܘa��5��E�*�d$=�̀���pž�<j�w���{=�u�?W&i�f����E*h\�l�nh��C.�/Z��ʺdc0	��9�E���Óf�)%<����G9=�y�s�*�9϶�:���{�ﷺc�V�1Ӣ�1��yT�=;K!��4b̪Q��O!�BkwZ����b͈�	{�-�t^�)�[C�?����������l�K�ݽ;�8"�U��Vn��q��&t��t,�檌Vw7S�Y"�yK��3��!��mB���-�����nv�J��H�7N03�*5;�*� �ʚ/ca���!_6�a��w}6T�f�ʋˇ�_��J��d������L������8�l�A��
6����h����h��R��^v�,�?��7|W���0e!ta3srʥ)��ȸb�����v�]I��[dk!��{#1n�MHՄ:`«,P��x�sr\4Md����9���w��I1��5
��0�z,G �"F1q&��L>�9�0`���a{'����x�8Nss�'���H߈ PZa7�V�����[	�/�,w�+��|����-�����r��1���Oj�����>���9F��(u������4h��3�QU-֖o3#������ZuD@�?\��N9x���b]��8��,/#'�eJ�9���g7�r$S�@;��s��K<qvǛ�f"D��m͐	V���4४����ѱ�ǋ�/v����x���$��䳮8vg+ݣu,�4g,w<h�V3y���u�=4�71��g����s�3μ���8���>�}��C����Crl�o�;e�~g��Aia�+&�zv�_luNL���N�����{����j� F�r��\]'Ȍ���[�p�7�>M�hr� hny(u(����&<���s�J`ğs��}���u�F�"stTF��ȟb{��Ѧ6h���m�c+ŢL�<f�8y$�Ƿ��� ��VvW��&��1�LС�o^�ѯ�%8G�h��?QZ���n^:$&�컛5�����z�>����~ӳ�K�wpf�V+��ئ�L[�z�!�j��G�p�����
�j���M���44W�9>���e�O3�K��XA��݈��DsO�l☃7q#�������f�䲲BE�1�o�|I~��p~�_��۵�W���w-cEc�*"�+�9�Ѳ��܉�s������P���d�7w}UW�x}����/n���w~ ���w炙�#0C��%3�^>��fL} 2*��깏�_���pe�X��|�
4�"3qT�Bi�\&H�i�����w$��s��&����e�n6�V�i���FSv��|*�ۭ��������eb����c|�p�J%H��d�ϯ�g@��;ލ���<����OM�������G�@�Jۑn����VL|\̞ �{?��O��!��y�����8����D)�~���'��k\�گ���>��3��J��vՈ՛7eTTn]�睻��$�_^<Ad�^7<@��K��ǋN@�so"�it\ñ'60m��P;���`��{{�i�!�H�;�e�L#��-]�kZ6��W��᝼Y[�����6Hr$��l=٬�z�[] }�"�_�іqc>������U��|Ζ�cȤ��R2�&S�n�b-;:4%�	y��[sz���aqQ�сiG(�����Vf>q�ed�����
d���۹o`�]E$8����ތ�� ���^�s[�񻷓�,�H�V`�Dd��$�c����Ɍ8ڥ��ވ˳��B����S(̤D-������U'��e������r,�}�(O>�n�m|{�Q$I9Dɏ�_��;@��7t{�^�ĺC;~�Q_Vt�\?�v�jNV�%C�:��h���w��xʶ���@\�/��Ơ�����з��z/��̾�Ȣ�੸1��m�<��!=$u�6:�d$Mr�O���7&޹�4��5��ƨJ���!g��7EN�m��\z�v�ǃ��;۱�N����u�������jp���WU�Q�s�]G9�N2Vx<t��z��p�l�ؕ5���c��\Mpn\<]�88y��JX�p.�e$:�-�U�;����KŞF8��;x1�uP7,���<Վ�u��'{��Q�w뭯L�:5nU��FѶ��<ז��P$ "�|��D��a!EA���n�Έ˞I�����[�:ɷE�8��U�î� 	2i6���E�V���Lg��� ����Fn�k�4�7#PB��/�<���	�7�<D��U�s&N�趷z �u�lO�0��0��ħ��m�"����t]�|�y=z�
T���(�L��=�B��b�lt�"�j������Bc�ȳ߾���~��^�x����v�B��҇u�q�H@���$;-� ��Î�m��o������Ɖn��oc��Vfa�@̒�E���Y�l�r9��_hx�	;�w���1ČN"ƣ��^7�<�Ps�F���Z��Ll.;Fj���[/����V�L�3O����ک��.�`�����rtb2�jvw��rt�>��ü| ��I�V|�!�E��X��kyt�H�%]��z�x����DE���W(H�LQD�m�c��F<�s�fv�O���ɟ��:3�\�4B�! ��Ϊ�g+2>���l�ø����{�躟d1 �BH-31��fc~#����.�9��"�v�ދ���}2J�m�����D]�	����k�Ír��%�l9 �'g�\�s@n��9�����~����5�qQ�DE�'����k�	���i�((�Ff=��w�p��~�?V���g�2wn�Gwt{��{�����j��f�{�F��=���������]�Q9�����G�3М-�yi�6KƬ��!�aFv)�7L��N��̚��gg/������͵��TP ��1�v-r��9n{��j�p���ﻜ:�g��2dF8Y�A��ݛ�*����̑tw2fO��Y�6=���p��;Ꟃ�&ey)$�	�+>���]�+�DkY�i��}�ͬM��L��0�wG7��5$@�&8"`�'�]BE�/>�5�zS����ݖCۃ�D�N�f�g���� PS���]�̙9�y�:���l
�w8E��툾��FXp�
5$�b��gވ�u�G�-ZS��j�2���ݻ��-���"l��ku�>���2�%�*���wX�hg1w�!��X�����ƋM$aݛꪻ}ݙ���X�'�x�d�fx�hB�xs�/3�o��Ww�ݞ���/l�d���O��@9��}���l]Q��xY����%2�`aυǽ��״q.?����ƉJ�������]�[ʻ�k�o*DQ4�o^nl���:�i'!r6�h�y��<���UB({޳u�_O�f6��v�(9^<k���r
r2�S�@+g�ͱ�o�z��u��wi�皏-�[\H��&T�$�i�:**�����0��v�7s5�l�����a�@̒�L/]��G\�ވ�Jv:�Q�{ks��x*��v�;�#���9��m��!���+}�}�)~Ʊu�V����	��(���"ٻ� ���kܝ\�����;י��lt��ڵ0X��R�rEw��?z�����fa2v:MQgY����=I+��e ~y�y�nͨ�h�{]4�i1{��L�|t�|a�߷�rL�p�͜��M��)��y_�N�.k(ϣvY�S'��F7�2��qtrYC�4��s��e(�;d��*�`���'1�h��w����g �:�Xv�޸ޞѻn�O�r'���1��.�+ݵ{��p�ްN�Z�b9�O;5��M����n9�b�"WvNq���^�R��{n�����1�ʆ�ء��Z:vc�l'Xw6nru��1^x���CËuI�4�V��U����ە8ݎ@IsX�+��绫�7�sR�j�W6�QPEh h��Yia�LI��F��bb!V�ʼp]u��ˮ�O'�����FC��5�ɥN8"A���'�c���ǻ���$g3� s{�5�8���D�
T6,K_W�P�|_p[��n�/s&t 6O���$�e�(&�;��{~9x��"�ݞ�C�=�5���r����(�P�����U�vɶ���wTƂ{���7[Ϗ}(" %!JI���ߣ�g\GD+P�՝ݿ]��iv�(rs�!2�h�dG-�p�ʖ�>�E�ݧ��ڊ.�J�Nn���Q�Ԉ2T�M�&8$�̸�������=C�Y���Ri#�Ғ$)!%@D5�vq�+>g�W�{��;s���^����V:���2���!t芔l��j
y�'3/e��S���C��Ű�iޔ3P���<��9�M��5�Y�n*��w����� �
+�@Y!�H,PA8ױ���a�L�l��75�8o�+e�	���6X��*7$7gz�Vd�����Ul�xt��{*���_�%��1�"���ވ���9�I����[��w/���|��8�H�-���-����T_���vѻY��̘�EW�$�&�i��p���)u(�y0��h��kc�+�jFl�r�C#���i'rF�a-��{ٙ߹Օ���?�|��N.����"Pd1v�բ��9t�,�v9%: fw�YR�I 1:�]��i2�g:�Кj�5��C�"���Zib{��H0{�P���s{Qӆ�k*X͍11W�z��v\ƵBV�O ��XcU���u��\�V����� ��~i5U�
�0����ύ�_�;��I(�#+�z ��IC�U\��~��}<p�_s��$)�0�hE�����ƨ��7W�~^ɉ}�$�P��0�9����P%�=����<�'v�t��q;n��GO�/3�����|�v/b��Ww}7����L��~���CتZ��}p��	$��b�>���:y �~�����Vg@�ϟz�D?�
m�3ǣ�cU.���:���������L�$(���7��d�9Օ����P_o��}�=�(!��5�[
�(�����[����Q2���wF���7��A&.�nn]j��+srg#E��l�,;�w���y�̏���z@F�A)R�]��n��^sG��O��|��<^ �B�E9d�ö.��
�ή�Ծ�^��ʠ>��b������5�-���eBCN���]�]uwn`��i.P�ժ�3ӻW�W6e/~g���\mS����U9�ҦJ������$eZ�����Unk۾��k�y�~$��z����"�	�v�z*�8ꊭ��ϗOb��������RIp�l�Ғb�;�uxn�4N^���T+��w�ނ�E�ÍFaaL���� 3��@��6X����_dZ�]Hl�Tޙ��w�m��R2�	�o��j�d��{�6�
,j�۰uE��"k�2����왫Fj��h{��xf��O<��ds
���>���S���߆+�-�ӏ�lp�D�<��M���y�W�zzr�|��U{{jӞ~�y3�coY��T;����.��z
��>+�6?a���Z�n�g���&=��.�3 #jĶ:�L'�/�Ψ����V�mt2f��&��`�����N`�:���#M����as�4N�f�w�/C��F��Bz�u��^�e��ɂ�Uq7C�wD�)�7��ĵ֙��A:�zk�G�Η�N~f��z/��|_�N�������K�b�`�ΌU����x�.pْ���Cѣ=QN'S+��;�o�����p���<8�Oo��s��q!����1����	�=��7	���Э1:Ne���$ğ!�:�;N��V*8eI>N{T8U���G=�'`O���g���� 7�Y�o�I�­��4%Q��,Mto���u��;��.�)�v����zp��qrE���F-{�N��[����Q�gT�U�n��Bae�U{��I��n����ne�Ѓ3Ε��J��u��Ño��ܼ��F�OV=����И�ק'�0{H���Y0���f�OX�p&�[$VL&4Ą�c�������u��d�q��Bɩ���������6M;=�<����E,]6�j�1�s-41S�N6��]���v��N74��� %�}��u"ͷ^x{��>��<��	�w��Ǻ2���u�C�P�ʁ;���d$��\o5�/N�nT^����rq�#չ�/;a�D	Ҝa�jV�y���^���:��,n.�WN�Iutq�-��:^m�^^;6�]�n��uu��7Kmq�R���u���ۺz��n]�š�<
�B�.1`� ^�n�� ��5��y{i�UȜ�	�iۑlC���Wg��8��*c��V���L[�{s�s��]:0��n��7'<�q���n{t�R��֖z���ǳ�v���Wk���r���+�P�^o��&��5�n��OI��/<�S�.����e�q���T�j}��2�=d�n�S���q�v��x�y��[���&1�N�Ǯ���؎��v�:��{F6��ܖ��7N��%<�=��}�<�Q	�i���<��`1!���c	��OI�˗�Q��;6���s��W��펝v*�Bj0S����X��*�c"�k�ss�g;�ŝ���-ή�hK���l����Nt��661�s��_k�8>���w��눻:0�kd3L�k�1�q�[�.69"u�kݒ��S')�v�v�+�[&\�t�my銷$;� 8�I�:��9���=��v.۞�:�`�N��ۉ,.�u�p3g���z�%;X�]�)W^2*v��c>�{/k���6��d՗�*V��n،�N����9{p�
���u��������u�n�����I���v��ە���X���{:�u�:�k���d8������ܸ���3R��Ռ�Gl��'��:���<�cn{8��A�"��LF��خ�y�sݍ]�^�����>�W��xa#�Q��u�ɝ���̯Dl1��W}�(���t�a���������x�0�	�1��ڮ1��Nײ��Y�D<�:֜h{>�8���u���w��<��gr�s�ƭcn ۜ�-�g����q��nμ,�m�qBp�v�1u�,v�n5�e�籼�v��ټu2m>$kkqq��#h�\�f�a[�����t�=sc/m]U�ڜsm��5���h��jd�;;Q�a2��fj+�)�fP���ٿ��%��]h���5y>w_�(sJIcj��9$�Y2g�4�N��K�$0r���l�Q`;�*{�:[���o�ڪ8�ǖh��[�{���L+C��Ղ/L��-�����N��O,�i��X�YPzpĨ;4q���i#��t������#gQx�[� �5����qy ���1}���p�j���h���.l0��V��2ސ��z�����]���\�5�,�-hF�t�0u�ws�W�>	����|�G�F���M���rd�����i�6�����n5�J3`dvi�1��-��ۈ���8p`F�;�(b�/)�.���P m����g�Hg<��+��Q��̢=�7!F�v׭U��V	ɾBr�{Y*�{���Ω��P���QY5��}�i[��>s]��dNc��^�R�-ᮧ��;�w�^h֓X��)x}�i�/�34������Z��._ ����L��}3F�2q�R�*a����V-� �T?E�˨��^~����z�4`�_x�1k��<��=�я��0�)����s Z:6p��R�nڙ�8tnd�++AeF`����y�{����A�r�u�kcť3�C�SIaZeu��Ӹ�a����:w|�*X̃6$�<��+�v��a��61h�[�9�G=��=�f�O�*Oq���J�za�,7���罉��04+�c��u�9�f���1�ґ�;(��:���Ӌ�;-���g�4 �?�7Ҟ����y�c)$fܚn@uz�{],q��@n��{M8$��3�t�G[��w]\4�[�	�W\P������*,�7[t���gsC3�ޞ;lr��C�Y�Wk�8�d��]quV�)��+^�k�L���a��\8⽖릳����9c�/�0�pt�l�?�,Q�1�cY��&U�Y������[��gh��V�w#�n�7u\t�)=-������͇1�c]����{/=;�����?`�?B������}�x�'!*B��99��ޞV*�Os�^�#����U���β�n�J�-�������]����l���c�8)2E��A��@��"w>��߄|tw���<�J7n@B�ԸN𷽪õ��}?Ey��G�-����%2�l������+v���{k��"�cɘk4�V��ݻ�@�j���t/�o���_~O� ���GXd|�JSJLY���O��䐫��ٴ��vE#F��[�%EQ�U�5L^
��vƫy;�={s�7��p�z2�cz��� v��F���ݛV�����r3���o<U�~~W�G6��oڻ�����'��;K�U��oàPɃx��\&�I�?������
��w���Y�y�������r�P@���
�2}}Wk��6��.�E��]٩w�W_��5$(��{��Y�H�:h�7g��X�Wk� �s̰�i76{ZPݥ�C>oh��xm�wC+� ����ӋOU��ː"�$�B$T���׾�^�y��̘���G}>Ŝ�} ��č��Z���>C��~�4�9��v���}йw�U7���q�"p��256bK�6������>��9�K4gͯ)�yzp�œ��+) �w8ܳ�2`���9���r�4r7$g��R�p#oR����\E���{8p�Rg_a�\�C{n�Ǽ+�Șr���a����;�f���Q���ھ�A'�4�eH�r�M�#Ra�|�E��5C�9�z�����s�(�Ǣ#��D��! ���nΎ�������n�Wkp[ٖ�lv���׬���E (\�8�j�����	����W�P��p�]����$�0[,)���z o�w�#۹�|�<�߽���#EHc�9�f/��j���.�j��z(M]�����K	<I�YM	(c�U�?,ɽ}�<Ip����<�z�z���3f�xv��f�nι���5.� u|�,Z��=%VJ9�}��N���T�e
��;���E[��]�Uv��־7�t|1b��Y0�1`.��s��9���)!d�	QTi��G9K��~1u}�n����t M����*������9���y��(�AvCۛ�z���q��ԄS�����Zo���Q\R���E�dw�ľ���Hi(D�bn���{�so���?����\#����Pl3�M�-ŋ>�^pCh���kMT�ت��bvN�d$`$Ƴ'hx�\S�ש.�ڊ�p�V�/ٞ|�I3	��_>ty�/C���.���|�ɉl�ٶs�qw��n��J5ӓ/�т��cE��0��w]ƌ�u[)E��v7+B5��ҝ�B2v��Z�<�9����J���ǵԝv�z׌q���q��s;K� ofJ�oP���e�a-�q��m�v�q��[���g�}bh�����~'����89JK�k��Ջ�ݳ�A�%pT�nϡc�Ӓ�w�rm�sf딏\uot���`���D]=���$�Ħ61���m�����s�m�� �V;d������5�mt�����'��{pFҙ�t+����|wϟ<��Ι�t�[�����n�:��湭�Y������Ha.���cb�v�`h�Fd�Ɔ�*8������jf��wO�p
��=�u�#���B��*DS�c�|���(����ėHmn=�Uy�s��,50�%����;J�h��� ��W�n��껙���8̑8Zpy3� I����krGER�G����͜bO�$˒$���d�<�����P��fM��^LIp��hVf�~l,d
( @��՜��#�A�L���7$[�x�|�GL�Mp�٭�(�2��#&@H��ã��.���q���� 7_W:3&w�O���0T�(��O�����G��T�����lS�M�7䚍�X���D��J��I�zZDd��
�O4�[�c�[d�0�_Q�����1h�{LX��f"10�b1�Zg8�緋���P�{E�$L���}��O{ާ��F�=��))�E"R@���z{W}5��E�f�+���ݎ9��˾q�MHcND�I�yϗU��
�޷��r��P���4�0Gn=r%��jG/[�9�:{z؍��X�)����ڦh�Z��P�mH2o�Xq�7s��:""�랕K��9Dʓ%%Q7s3�;��/-�h}�^������yBQ2T�((D�!��������0l�g}��&*>�9t�1�ky��~���x��ds^.�t7�<�ή�Ӷ�����M�Tb�>�^�v�_+�)Ǳ���A"J"�H�� ��D;�kʹ�Ck^��$MRjYq����Όɼ�"^���ER���A���@�����8ݞ�p�w��.��e��x>���NCa��痞�URcwb��۟]Uq�s�N��+B�-�l݆`cNH�)�`!� A2�j_>���./�-�ǟz�̽��^LK�����P)�*dE����#��띞�����53e�����<��B$S�' ǝ>���>q�΁A��_k���}�;��X2J
 �2�2�G���8�⃜q+k�Srat�:�*M�:aevF�3�	Ơg[�"���{�X�rѨ�1.{V�8��*�0Q�}�m.�r����HFڋ�V��/3L.{�3�`�����=�~]}�8H$��� � ��� �$RJ�[�v��'`1�q8Z($Q�s3�	���#��M_9�~��sǶ�/�@�M�	b�aJ�:$���ݎ�)��yX�4�Q� �5��07Pn@܍$�I%1t[����w};׳ []!���䌎Ti�d-�Y߼׆g�U��{��������j������'ЂF1-�>���LIp�PG�?�_~�^���H�i�����o�}w];�F�Hڥ��g˸�Ľ�װ�"Q�$n9#1}��W�(s���Ncz�L�li����Mt�x,��!ǯs6������<�7�y�`��>�5i�-��f��%p��/.������iZ��U=v!�1�	��Xk�n�n��:�
���qpl��mX�v��`�i������w��c�y�{��Ń��s����B��&�i��������x������Cۓ��7lv_2��gM�m�f�/����'3�vǞ!os�敢{�������U����}S�ܧ���>Nz�3=��Ώ\d�m:+�բy�� p8|]t����3�7�����}vy�D{f)/Uk�*$P$�Q��	m�:�)�V�������n,e��b�O=A��:�Q�9��WZ��ѧV���=�9�#j���6�ftG�z!#l��}��>��B�P�Bm��>C���[��s7��������_D���A@IAn7�4�R�"#��f1����:)	L�I2$����ފ��UN��DL��KCL W��H��5=�b����L=�������OxP��)x�K��,��2��͹��ݜ�c���d�b�[n����E�]]*`ʙ� ���Ec��舊�{�[�~/S��K@P!�o9�{G��m����>&��fFq�]u�z���|%�/�e;}�쟮t�,6i;?_�ހ�Ԭ����*�mu;���v�s�R���\�+w��E�C���$Y�#�#N{lI���w�\�U��$�ߩHf@��o��;��*�"!�ޚ����:�1��A)M��P�{3z��d������Y����M�H�a�ZQE�z���<���ބ��ꭏA����F�7Zw�;�GX.��X3ϻp���:�����X�j烁+ ̷	Z��($V���MU�5S};~�DFe&cz��2X��H�R ��̢R��ν��7w��{����m>ڠ��p5�dr�L!#Ra�y{�2jr���-��ub]v0�nPp*�nF�P,X�ץ�\껚�sv�d1/eo�v�H�sWTy�F�/~s�c��D��^�����y�n,�l�Q��c/��N+)y񓠣��^��8B�1tG|=�������)=s�FN)۽������s{�nTed�f�}�i"�g�.OF#�9�\|���)�C���x�w&�n��L^��{��цz[q=W��W�����C٬zc6G]�w����h^���{Ů��;�&��#YV�P�SM��V!�'X�}=brl��;�G�������yr���x�K���mf<�3ޞ}�$�n,��^�I�|K�<��d~SsF�;�{<���ʄ{��lK&�vc&�Uo�̝3*�r#{���틹�3U��Ϗ$!Z�����ZA�o�^�S�NTU`L���d;��ރ���������Y��GJ���ո���f��fgz�!�������{g`�;��*�^ʩ��Y��(���[�±W*�]<
��1�܃4]J��:;���ϐ����+dv[�-�ޮ��@�V+Ls��v��Q���ٜ,T�w��h�.w`���:��ߒp��}�Fܝ����Pv�����M�$!�Z���˧+o:�a6e�gZ����y���vW-kDF�^��Oܔ�2~���D��In��U�謻R��ej���~(��,c�~���	��,�`{�z�J��y�rDV�U3�5v�'��Tλ��5A��k�������W'��/��U�{�a�@�������g��7xu���7�.N���3B�m�u�(�(EfU�t'�n�9�W�<�����2," L�Ȗ5�+BN2�h����x�n�n��]Q�V�� 4���}��AD��d�/P�`���0D
^�d�w���l�ƭB��AK����cj����k>q �o���q���,�!�D���霯 ;������p#�(P�����kS`�&��Y�X�>7�ό� V02��Ǻ��ۃ�X�t��!ɥ��Z�iL�(P��4���3pX�&m�[7П�z��G�-�2S�x�D�A�0���[F�������E�����=.{���{�&�,�g\���|Z'_�p�q�p�d|6A˰�����坷��3�伮2�)��ᚎ������_����S�q`{������*�7�B���͡����ԇ��ZN2�G�������+����9�յ�ۤQ�F������ o�gaǂ�M�Jx�� o���C�9�u�T��I���Db��rz�7ϝ��W���H�� 4��Fxn,	��;�t��c
��Lj�9�I"x熜�{��6I�����5.�����FRo�����]8}�{�fŕaK�'�� Fى����5x�.�3��{�cl�Ň�ܽ\;./n�צzǱX���Y��9�κ\B��ڎ�����`�c�<�����^:��K���+]�Lo��Z4ڔ�+�1�H+�!�{p>^�mJPa�<eP��0;-!�ן`_" J!�@��R4v<�Vg��I�;�0&J@E	$ī����֛m>��w���� ��ݭ��z�.��6�h)����]����f}��y�y˄��w��gІ�N��"�a����������-��gVz)��u�ϫM$��F���7q�vc��z=2�Uh�y�̆9$H�����n�j��r�t�/�wʪ���e(��k�r�7���bz"4{�1=��}QU?N�.H�h�\%�s&z��ê��;�����fG[�=����^��\/� i��ʻGMF|�&�La����};��\ջt���}[7q-kܝ9�o�-�M���t��f}�m���D��M"��c,�)�E	��������KH�l$����wڪ���3��&$�qI�@`��d���0X0�W]��k�_t�r+3Į��V���#sb��,��z!Ge�����Ũ}�v���>O3�p]�;=�8�Q%&3��'����3�;��s�Y��O��^�)����e�ĸ�Ү�߅��P��83��&%��G��da��
{��o��3�r�GQ�Ns���aI&aA)RA�>�M��� ��:;{5%�ԕ<5S=vw����2����UZ�)qqa�9�{�^��fv��AyC��-j*���r��t�+��g�yoM� K0��_^4��s=��Hófj
����:#E��	7mk��Ol;�g-�f�v�����u��Q�r��S/n$Iv+
��n��u����n��G��]@b�����˲0���]d_�ݼ�;�Vt��s�̢n.;S�	��v�3Ӽ�ac=q�;s���⃫�v�ʉ����m�ֺ����7lĖ��#�W`�u>�Χ���"63��^��6��;v#�<I\��||���^�~�#lE%�~�PDWF�y��aT�Z �؂�S�`�����r[7-�/֐�m=q����-
� �و����\��Z����<��ޏ]�ީS��OI��JL$
AV��;^�A��f�{��~����q�&[��!%(����@D�n�oERǴ��E ��w�0���{9#IG!��&�)Mi���}������X�;U]]�̍��ҙl�ȌN�Q�e}֪���c���fj��b�wg}�C�|~@��u\θ�n�2`��Y��Ke����0���l�V�ۊy�V;"�������ɷ��˫���b?��wb��rf7�N���F[j)ak��q�;���-�/>t&�ޛܚ��v:�^D����wy^~:v��r�ރ��u�B���pXª�U�U�#=5�������w2f�c�*<H�������c'{*��F�|" ����	����
ŀ���{�:�ֳ�M�m���M��}�/km��FF��$RR�#�}��c\�L�6E��w{>j������fV����s�����e�%Gڪ{�1���E��A?K��Ö��m�c}�:v�u���m�
qt�R먈���J:�{Nwnw�֪�em�ֺ�˚wWi�ȑK�H���I)'M���R9�����n��0�Z�\�v�ǜp�!
8�M�sb�����l��{�Vf��WG��s���C� �I@Ll���>�L����p���ў/�D_M/<�z)+ʀY;�+K ����L��\Y�s8&u�n�S	�ک��Fu�{W\_ϵw����x���5����X#$�Q��$@\�Wm��pmn�+���(D��Rvw��n����<t�����C��N���!!!#��fT�z"7wsْ���&[�����{g���-V��K��W9���8�7���45�4�:m�/Q�իv�a�1Iڒ,IL������wgN�ڻ&\oDG�]�Ү�~�ϱ4$@�2`iI[�g�\�{ފʩ��9Y����j�3r.�=���lL���<M�_cۭ���RW���B﷟�X�TuͫJV�vJJQJ6\��{{��s+2\ߞ#�2zysafg�5.���.��~K��(t6�J�����/zt�8�u�dv���6��W^�Ly�&��t������v��ݦ�=���ϯ��.������Q���@���w�9�%�Z"@ԓvO���?6���Q�I�g~ﲳ!�$�E|E}��&H"$ �d�S�nDp�g�Rn�w'W,���x����F��L����~�Wd�v:��-3���7w~��n�����h"����e�f'������|9u${�831��s�Pݓޝ#�8#���R0�׻����9ͭހ!�Pzɢe�oefo��I�����Q@�̞�S��ѻ����&ck��'j����]��V:[�ېFDm��Z�ܷi�B}���&j�;��b�َ�"��?Ne�t\����,�OD�WM�jV`u�rD�iP�m^'s;���_OM�[l���l�oCޞ�Kg4����t�Q�0���z�����8��ų��t����&�F���Q���k���غ\�9N��2��B���R�;��O/��25m��e��r��9!�4D�[;����c�[͹8ޟ'�m�E��j�۲�&���nӋ�ݻ�ݶ��t�� �,4�a�n\�Bûvۗ��tj�N�k'N��s��n�2��5q]lr�k�P�9��k�k�ĝ\�霽�	q6�-�'E� �Z�Z�M�v��m�r�ϯ������wqHӺN[��Ę��S�g]��u�R�rv����e�Bn@�00с�c-'�ZY����35D���{�Cmi�Tf��BEN@�	6n����(eϾ�љ���w�m|9{��v��qB��(�m6�Y���|3٘Y�T~"=K΍����{8#���7m�ߨQ]��	ion��2�l{л�7dO��$�P ��Q��7���vn�M
�����f3��0e�}�g;��)�J%T���q�n��n���}s=���y�vf�x�k�\�P����	����㘏o�ݖt+]��>~�����\-0�,)"z����U���'�_j���M]z�W9��@�ΰ�S^Mt����=L�~�5��xwj��fa�̧ܫo;�q�s>f8:ɸ0�  �@i��W���v7���.i#BwO�}x���wy><�6��<�@�Q�L�FVi[z�>�����_���ۋ�?8�I0(��*
�_G�;f��;�K�����=
5p�J�[�<�ϣR6�dFě7}˫�?{�o�Ff;��VL��5]�Ѣ��	��b$r�������f�"і�n�0u��ΝW���g��?�����ؿ]�gB��'���z!�uz����	,�Ț��h����x�� fȸ;n��7h��~��b}tA����Ա�?�f�yuwr��Pߔ��h��|lC��4�Jf�{T]���̜�k2ֈ�oi�p���e�Y�۹����/��EhIZ������F��f�zv_�l�I��H"�)"�v�w\Mˑr�9�b���B4�>��2���	x�;8z[PIM#$A��w�Ur�<�c�:r�0��T�t{�5�o5��O�$�@��JRHɕ�-𸻳���'xvB�iJ�j�_��6r�.�!G����"�X�i�d������=�p����nǳɲ&PH�I�� ���}P�l�H�=Y[����
�ݾq�6�zz�	p��$-YxA���=
�V�7�q빓�X��{B���=ߊϠr7%&�m �u������l܋���e�i�c�1�>��т�16�R<y�;�r���F2��4s�ܓ���x'�'�d�G�q1��i��u��\�����[}��I�Z5E3o*k�����U޸�T����N����1Q����k�KF��3_��]��]��A	!˜�7uȒI^������an(�DƎ; ������G�W�G�6l�"�֭w{���߰ʧ[zf��XXl�ݩCt�[ۊ�뎮��ؔ��6|�t3���q���v{%K�����+1:����܏���ee�蛛$�n��E�&�kݟ_g^��_�޳�n�'b����gj�f�<p(1*�����=��Q�0�Y}�_C:E����ǻ6�yȚ:��c`���7� ���ӳ$���m�Ϯ�����rV����)P)(�T%�M͓��F<�c w���NN���sc�i�j�����~�����Li! �I���������mU��ݭ�[j��mV�� @'�H (�H!o�C;��$?@ /����������۟���?�������?a���O��|������g�����I'��������o���B$�rB$����x~a�O��~����?�H@$�?�G��?�����_�p�K���w6��mil���m��ii[6�Y��J���&ڋl֛jŶY���i�jZj�kM�mi��֚�mimf֚�mikf�m�6���kJ�Vҭ�ZV�kJ�U5�kM�6��f֚���jʴ�ҪmikKT���6���Z[SkJ���Օ���kJ���֛ZU�֖�֚���U�Zm�m�Vͭ-��Ҷͭ6�miVͭ*�ڕ��KZV�kM�-�mi[M�6�j�m���[M�5��Zj�j�[T�SU��MmR�-kMl�U6���mi�����Kl�k6Ե��R�ֲͬ��ʴ��)��j�6�M����-��mik*�֖�V�UM�*ٵ���jmjZ�Z�ZkT��j�kMm�֚�����[R�ٵ��ٵ��ͭ5m6��Y���R���6��m6��i���ͭ-jZ�mSkKV�Z[m6��ZmiV�kM��֖��ZV�miZ�j���Z[m�m5m�kKZ��ҭZkR�ږ��ڦ֚�i��ڪmikZ�Zj�M�6�eZkmJ���J�Uf�����[i���KZj�V�m+R�M��M�*���j�Z[l��kf֕�����ZҫRږ�M�+[M�+m�ږ��l�Z�T�ڦ�5���-[f֕��֕m5ikR�-T��mM�6����kM�miU6�ڛim���6��5iT����Y��j�R�e5Jk)���5)���5��f�m)iMR����֚�ZYZ�6��6���ZV�֚�mi�f֕Y��֚�mJ�[f֕e��6�����kM�֛M�56��Zi�J�Zf֖mie�6ZҚ��ZY��kjSkI����mi�ٛY�֖mM-S5�6��m4��6��kM6���-i6��֙mi6�mRm���������-�%)L�[d��-�6��ZM�)��Z�[fmi��)���)j����Ze�3ZJl��M�%��V�ͭZf�&�5JlS)e%��)R��ckI���ѵ�V�ե-�5h�Q��U�kEmImi6�����&֓kI��Z�m�J��m�Z-U?��魭��V��MUI��V�TUh��-�)5�mkZ�Z�h�1IU���(֊�5kM�jj�jU-f�mI�J��M�)��mM-��YM�*m�SmJ[jM�6mS*��S6�͵3mJU�6�M�&ړmJm���3Z�j��IkKJ�f֔ID�c8�F�?���#�d�I"~'Ǻ��q�~��~@$�~����������L7���?I�������	$��������~�M��<��	$��H@$�I�"oP$I'��F���	$�����3�l��G�L�+%$ I?������9! �I�4~S5�~���������1$ I??���! �I��_u)O����1�,����?��+���M�w$ I/K��&�����O��p���I'�)��M\��I$��?��������?��LPVI��Y�11��7�@��Ϲ�d/���+G��          x}P@  ���"��  �@  ��E+p ��q�zYh�F�v;r��֍�us�5���J��wn��{�6��]�Ӗ����}�:{������)| �����gF�Ֆ3��KF��ʵ�^:��'ªT����_�&�5��+�*�� �#�y���B��[v�mi�IHӲ>�;�62�7�z��v�w���M��v�Mv��}�J_  1�������m�m���[os����=k�T��X��^��q��Ӧ��ݏ�G�: ��nU�=h�K��O����מּ��3l|kh������㻔�Z���h    S� �J�� 	��  1�LIJ�       �ʨ��        ���T��@     �IT M 4  @B I�M ��i=�=54f�i��O)侑�@$��I AB@�$.䄐 y!���BT!$���������)���Iб�!!VL�jC�� H���� ,�5��L?/�/� �t/�~�Rt��X}����?c�?bs��h����CܑNd��s6ɼ����L@3K����nܹie/eݙWk��#&v�`�]�AW�&�&�Z��\�*��F��!g4wGk�;�ް���V���c�wc��Q�o7�[�{pq��p��SN�5�;u�(�O73��75��N��qˀ�4�O��8�:s,dzg.ܙm$k]'w\�C� ]���id:s����nh��U$��u+;�����֭ؗiHR�4ɛ0�Ï��^/nSw
�R���ݬq�`�_GHӽw�5�v.fˇRC^��$�޷q`ː��sz�#i*�fmւ ���ڒ�z�
��Q�Z4ʉ����x����r/�i͎<��MP^;�5�%���$���:���Rq5���h����m�엶)(G�b����G����1�r�x�K'*���X��.W��2�3�e����L1f�;F�.iTSlu�*+�!\�����Ɉ;[Y����Qe�F>K1��i�K`Y��Xp)�G%T&tS�A˨p �ݛ���]y+\�Eõ�Z���gj�P]�n7&���������Mx�#��OU�d�]�2f��ݚ(���#�\��(��:h*�p޴6
Q
���t;MOb��(���mٯ��q�ʐhww7��XJFx7��Zn�>߅�~��2c
`�gn+2
�tu����ƕ�6pZn�dE	7_��Q9�U�[��q�q�A����u<*%�7!'TX���͆	��r��k�a(nˣr�rنS���쉝�i�8r�*9��){�1'�h�o8\�4�Z�.�yU�M�m}��=���`���Q<h�����z�V���>�)�I�X�N��`)��5F��e�ˈ"��:�#3D�6MH�s��/ۺ����A5A�=�XN�no�қ�8,f�BuF��.����{d�4��p7L6��'L��L�Uf5��4;b1>tO i�;&��Ꝇт���e��'�'iİ��2�E�:dі8L';�Ѩ�3r�4E�F�RԺ3Ϋ���q�:B�:��ˤ�n���$y���U�.¯ �#�-�M��i2Mdn���Gb��f�8�y^��f��x �UO���:Y�ַR���=���@����q��� lC�F#j�:5�U���\�㳙�n!�i�gfvoU��F�%�n��éE�f<��$k\��K�l��>�,ڮi�9	�h�D�(|C���"7���gu�%E�[g�u;`a޺�i�`Q����ȟ�yHQk��&A�����4��*v�C"�ݧ�O��p쵫�.7�!��8+����m�>�/������]u�r��6����Ȁ����Gs�j�U���N�Ulcꃎ�]5���.n��*��-&$٤� �(ɫ����V��kƞ

�j坻2�0E���p�a�����Z�R,-��^OX3{�r��V���l�1��%4m��h�]��z7j��;w���Nb0Du"�c�x��&�#�˂C�xp��V��#�8�i���4*�� �$vʡx.Y"]$����a�]�;���ueѺ��S��Ew�6L�W_�CN��ٮ��ir���5`.i��U�a�]�e�����V�C�x�V�'��{�f'��w%Z�n�� ��o��&�{okA�;�Isuʕ��IC
�����c��ƎڤմS�^n'^��Y{�
��n���n fAzө&ɍ[���4�q�:_(���sU����A��G^˪�Yn<���L��tAk�V#J�gg8^-�ݭ+��L���#ʶ��qm}r�0�=e'~QG�AWv����1�}&i�:��h�构��6���̵!�Ѥ�e�����5��p>�v��N+�Ŋ��8�ޘ�W�.��|h�Y�,7;A��
H�b|��y�v`�X8h�G���%���A8�,b	Y��`Me��]�#-���;�����ABX�3jV�T�5��]��Z���]�)��hڠS���B�ܜwy�.�;Ax�`��������0$��y.w^�l�(֥}�c>��o֡_(�<��8F%��V��j(L3t]Y�{q��y�������	Ww���yy�t}���G�?���C'�E���8��(��>'�|��:>Xt䲬�ܺ�Ͷ��v�q^ܜ�;��l2����^ٻ%�9o"ݓ��v���������Żl�g��s�;�rq��Ĉ���,�&H��"��M�[NT۱9����[���Xw� &�A�l��ሕG[�e�;<t돻�G�S�>�{DbB�;�S��bǺ�d�N�ϭ��Z���̀�����n�Q�t��b9���w��v��������:A�+�wU���F����'gtK �V;q�"s�z��dbh�<�mQR&s0ٟ�� 6��6w,k���~�l�A�v-�uہn�l]�O��,Ӵ�ݹݱ���^������v㢟\ݹ9����nl]��m���wK�"=ngm�r4A��R8Ԫ�SExoA��ۈ��)g ^5��n�q���qm�H�L����d*o��0]���C�/oڹ��<6��;b�C��q̣�:��1Z�k�+����q.��`ȷ8k�kӃe�t�3���1]���m8���n:�q]���Kێ���m��=��`�9�э��B�n��t�7Q����.�&��CS��o5�W�(��3+*��&[��i�M�r��y��6��z��.�˸�[�ֶM�9"z!�6w\x��r�P�n��)��K�m��5��m�F��G���Prl�����J�7q�@l�a�zݱ�Z8��z�(�k���h�Q��z#`簪����x3g\[3���lێ�e��v_=r96u��l���x;�?9�{rY��Zr�3�ٮ4{�Aڈ�����n�,�H��,m[;����۝-�qݚ�o��σ�N���8r�2���r�qd��>D&���℔�n�,�lY�1u�;^T3���uu��C��/�N~{v�n���8�\�����pog(��ؾ|��7���X��+�ۋ;؜�|v6�2lN8�o41r�p�P@�1��z�n�;d�1�zS��ϱi�"<���f�x��n�WK"�M��U5JY(�+�ܹ˲StW12���/V�5�mѰ����jG��vCF�]z,{.��ɕ�f���٦�̓*�Y��@�Ev��6'��lT�.��ʞv��vpP��=m���[����Q3m�*J�N#�9������L�Ȼ���F0:m�)v�;��բ����NTco�º�t{�������uۘh����]g����t�X���Y�|��'l��m��f�-w��?jH���trBVԚ�F��E&2�q(�BR��5����L����{u�V�Ө�;S:몵�h���%�ˊ�����q�
wROr�w��>0��y�쭱����Kts&��WYgs�mל�Zy�Q���o�*�[ǀ��@d���5r9�n�hT��ktg��zѷ�h5������EE%N�U�� �c����`�d��YK-v�p�뉩��z�z��QnMk/U�7-��mV�m�Vr���5p�ɑے�^fg�je�u~߇ϟ	⣈b���^j����u�b��^�g[�Qh��:WO�vE/]����Omz���P�Ԍܬ�n.U��\�oNw\��Ԫt�yݎ�+Fb4�`��닸�k�g�����]�]+��8�p�H`>��� @�?�T 1J��~��ܩ_
�s����K����x��1�|�jk�91W{r��p�ވc�B�笑��ym�:u�䊧m�G�Е�������m����u�~Ȱ�Zf�f���/m�4��9צ���n���U���Z�t^�[Y=�������d������};=�s�Bz���#�]���V��uwh܏��{�kʾ[ 0U�E��#E?�����;�^���e�P�=���@=F���{(}����k�)��3o�����#rf4�����>Gn�g69���ہQ���x�W'�q�%��̤���#�$Vg����Z]�}��g���a��h��zo�'��a��r�P��!���Cnzד6��ז�9��f5����D�>E6�^�w���}w|v�,�1C��:������L�}y�sZ�rr�,y}���>S���5�ô��OB��'7�ZU����r����˶��ڽ� ��D��ٸ�����z.�%8i@�����Ia�t{կ=��>�&j��ǒ�ѣO�8,�o{��h����}�����;�G��]��Q =����{~�įv�늼-��P��/�٦�~���G,�e�D�zȳm^�V��x�Fߛ�yWQ�:��y�䟩��5'�ûQ۠
�����,�Y��3`�YB6.F��ƙʜR��-ӛ�컍�+
I	���:��8��}�{���#�N��4�j���Y��t"����j�Rb�kP�9����������9amh��8�ؐ���`�ã�#�A���|�n�c��r���9��>�ZY���͖�\�9^6.;_����;�I���yh]�'�SR��%�y�'g��v�+�N�L�����N#��m쇎p<r0{tsɸN�ӕ��ss�k`��=Ч���b������,�;�y��V���˛���ǒu�-�}�����3Q���.������7��"Y�xS���j�����{s�x�6[�f�`�yūwn���^�^$b�m�OΩ|��}pH4��'����i�W%d�y0F��K�����{�Vۈn�6x [�����w���8��V|�NW�l$2��z�h^�Ԗ>���=���ޕ�p�c�6�
���K�U�'	އ�{nB"�=�A�]��2��7�~�=�D�����7N
_w��׾�l�}�s�^�vN��b��u�|u���N�G佹Wl+������=$ޘ��V횳�ȫ+ׯ����� �h� ���kؠc���L�� �C���7U6�~S��^�z�^�,5{o������{V��ս���K��I�ooM�M���#j/-��u��ǳn�ӏ	
���s��;�o{7Hڽ0�����
ٹ�� 3}�n$�Ӛ��N4�=�}����YOF5����ݓ6I�l�@����)���nL��٢{�ܝ�R��<ke�����FW7g�ss���#���4��3e�=C��J�H��r�=��Ӈ��u{d�>��aݩ�|��/�F�tq��ǾG�Jƞl
-m�Bkm-�ǁ���hn
.��"G�qh��\�Zv�D����5��$g�ؔݩ�;}��t��˘
��'�1�9z����'\ya�hk ��G����\�?|�@�sw@~*!�1C����w��^�X��Zb�3� $��D)�f�g�cyG�ޞ͍�/yo�g|,������l�T�Lwįl4_{o�@b$-�f�P�2�&Ћ��K>^É,������-�,�v�ۧ^��s=I1��=�nE�=�n����1���U�Nm�{*�r��4!�6zٿ?�/�h�FQ�l����s�`;#B�k�nn'��N��=X1�x�s�����"�e��;���3�a���׮�{�سÌ{0��3{vk���Z%��ڕk-ڱF��8�֌9B2�Eg�|r���B��^,Cb�ުc^�f�Of�O&�zʥ�i�7��'v�k�n�ӯȅ9���w$�����~W��kalVZ��wm�x���J�}��=�,}>{���2{L����-=��Eޱg�E�_R�6:f&rvb2�B�8 �[��M���ᑷ��妎 _B��4����? � `���H�E��[f�/b;W��{��=��ގ�<���F����������SN*��f37F��R��lm�ݶ�uNs��(�:u��"���8{�q�S[^�F�xܻZ�.:�0���{��4�ld��1�q�����XݯYڈ�Lxڶ���v8.�����\�x�&�7+>=s���׎b<�Zn���9Wi�����kc	�hA��rx�x�Nwi��ڋ=�v���p:��\������@;���u����q	q�Kv�Mܵ�nG���xZq��3�eyW����4���6�n,�ɳs��l�;����zձ�ys��rW=���Z�IZ5��O?��}����<�W�a�"3z>�L�-�0��1�HcP/s<�?n�����k����ͷ�&��(���ъ��A5����g"{��4㗏a�r-�U���觸1��b�NW.�ՕW���������Q��e_(��(L��	�[ҵ��{4矽��x�q�m��x�3ң�S;�}� |*4������V���|��<7x�����_<X� ����$�jo&0��=[T�dV���y�i�����ه��ه�uu�n����)��C��L���m�mu�"�݋�˞s@�DX
*AX���(3�F�2�\��q�܈���ja����f|�0�����A�A��f]�1�"��Z"���S�m�6�b5�V>�����Q[�W Z�v�"����O��~ٞC�-��:���V�FOf���F�z���Ǽ���\�j�
�H������l�PD�+ӏ��w6ɍ�T����O���RC'�n���;��qAu�Ռ�٥
9pݮPM �I�e��-n�$�$f�H�q���:m�a^)2�����?u�i
����J���,��wsM1t�?Y4�:Ö�����	�ؠ��B�TTU��UYZ��k�{��[�x��\�4� h8%4D99�|�C������n�uߋ�������I�4>����Qވ*t����.ӡϠ�`�j+#�N��х+;��J7<�ۊ�{])q��0��	'�e|J�X�V���=��+����o����4g�Q͹��֮�_�����<"+O7ft� �n��K��L38�f��r���n3�UKH��S��#�}�Ye�n��n��71�U�Q�@�w:y��}SY2pi���Kdq����l��B����3���n;p(�״'5����f�es��T��Z�n�ߣ��X�Ĩ��UA]�5s�t�Ƞ8Y@+��lw�t��x���ʙf}��rcU�_��ih|6���n�'��m}QO
������v_V���#����K+���>�7g*�T'�����νI�1�syَ��s�9�E������Jь�	�e���w�Js5��o�|�X�;�����v��9�0�u�;c�+crڛ|��f�95s�gp}k2 t�Gfvcu������=s$�F]�U�M����Y$�+P�h*V[U֕mE-�AAq���G��2v>���{߷����i��%���V�),be��	�-�@�,��q8H���ҟ��S,ȓ1��7z$"�?k��X�y1%h�+K�jcD�sǒ��+s�t~H�e��l�����:��x�D�^���.����F�,t����N�,ѪqqA8����ծsڨ�܃�G��8&�*�ʩ}�o���Ш��8��Ȯ�f*��U�i�չ�ܺ���8�ݥ��6�YGYX=J��L����q0�a���*�� mA���X&�7�3�!`�uZyI��G�A�4B�ؖ�+-�F"n軼�уW*i�.&j�X��!�߾�(��;���N�!��������O!_ej\>��Q�/�&:ֶ����P�C���+\�m����TD�|��w�r�TͺT�DX�֘@�C��5����Uƨ �_
��X�
�cm�Q5�3��F��q�����,�@l����yHE�}�W׹X"���d�R��є�RXm�s�wc�Q�yFU��c#�f��kϿf���ý.t|�>='f�s�QEbèD�`���ٻ�!!�/�������n��g �_�������������!�a`}z�"��]�o�w��yIQw+vsl�*v�&��'&��8��sN8��Nuiy�������M��c6d�װ����E"{=_@���.k|�<��b�f�Cu�-��mFK+��q]4;�8a�T����b�'8��q�~T���<�Y���槬gw�=���~ �d�O|x�ƅ�&�2��Hu/�l�kB� >�e�t�,��+�x��=��n/a'{�A��Uh W�
�B2Nf��U�ݺ2ti�vݿ��%$��s����O��f{���1cy4|��x���-g~<�c�=�A�%Fz=�����fL���@�L��H�y��om�x�ݪh��*�Y��M�;u󅭃��Fc�0]C�8�Լ�م#&�}����d�AA*,Lm�����"�l*���n��ʏ�]���A�P׷�K���W�]{�u�����6�򅀅�z��J%f�ѓ�c�%4���i1�ǧ�e���}o2g̼M�2��
8�=m�VR��NN�$fS���ص.{s��j��\��0i�2�=�+h�*
VF�U�e�k���/Z��=��N<%�<d�.]$!*��E(�a%I��9t��ކ�������U�Y�p@co̜���/Y�n\�`��� S��{{瞧�A�3��5�vf�?eֻPV����f�1&�i]�����z��A�BҖ"��h��͸�g�qn&�<;G5��]՜�[�ݽ�ö{�6 �Z���.H쫻��j���hh���f�߽��8򈠰m��m��
kzm�\�ik+r�#�O$�3�ʙ'��o��ƾ]I�~��n��3١ci�&9\4���s���CG*�e�緭Uޖ�H��.���X��.�c:��L{�����̽�A�{�ӏ�u��E��\|���L����X��1�,boG5�u�k3綪<��ǭ\�<����R�;�%��Z#D[e��}r��ޮ��8w�9�׌M#	%���=o���m!z����q�"p�����n�>��/�/���/g�Jy²�l+����Z��+�y?_E|brV�^*�=[F��H�����5��F�ک�QI�w�a�<�α���g9�����Ԭ"!Z��lO���b����T�6�^!�Uf��Ws����<��J�g^�@~�׫���"��E�5�a)r;����q�@�Ƿ��l����m+���}������Y&�7��b�AX����cƨ������/R1������#u!�kv�q�c�� _	�c<	��������EĄL�:�Ŝ,���s̒���NX��K
��gݫ����$�_&��-���\ko�ھj��I^=����0��,�F_a�޶:ц�	W97�^��HA�F��I����L >����.�<!6=[{!���T	�م�����M'�W�U2���\ܼ�ֹ2��|��/X��v��]��GBm뵄�u�:pk���U��گ~�=����}�5�f�4�Q�R!U@��a,A�3�щJE����4|�+[�x��%�@�p�65X���}�^e�&�R��E�ԏ���UTLl[H��śq�M%�+3�b�S�{����G{γ�-y��c�:<�HTܯIc9�͞��_aaaZ߽�L��]�j��t����:8�ȧ���_��EF<�EX} {�3��ߧRW��=f����n���D߷~�*�+=
@)뛑ԘKH��1�OX���,�c	`��jE�j��܄�nI[nK�,��)T�z�[3{�O=�x�����
�zW����k�*`�2���ړq��fꋺ���B˳�{0(���[U�@����í����
�܎�,T�Uw�{�2����Ж�����CV{�%�
��U�V�:���7�+�(�w��$7��z��~�n�t�:������	)r��cr<Ch�u����^�U{�*���i�g���ˏ��#c�dr�Ѯ����b�QQVC���fW�}o���19�����__��$TN:�p���R��abܻnYE��� �%���~��p�Y,�aMf�w9�S���B<ⶶ�7˜��^��u�ei)�MI�T��(���O�� �y-4 ̚�T������S�T��|>��%Ǯ�	3U=��Dn���p��Ҩ�n�_�SS�C�<���Z��v�ÿwx�F3��������Cg���g� r9��6�"��R���d��u�eF��%��&�6����w��x�z�n��򵫑ХPAt\n��S}ɺ�Q`���N:��u	]�J�7��N�r�Ӹ�Ǥ��{F����z�یbt���eLT�OMH0��<���H�R�%����Z�-�Я����PA<0�� >'tf�Mm�k]����O@��;l_]!e���R=�oF��d¥˥�zfr�v�ͷ`����n�]jE�ǮD�K��g��q�9�[�K���v��[�3nύt�.�pl����d��� �ǭ�z�a�c�^s����@u�Fك>�M��+�諃�����˛�d�q��N(Hv��M�v���D�^���;�@N�v3ўb�x˱n�j���b7m��]����8^���=qۃ�d�^r�8���h�����k1�v�̗WF���]"3f��+��c7OD�K�©d�Id�WW��Z��xs�i�~���Q�vh`1����8����_I�$j{�K�۱P<闯�L���R:w�<�6�v�VxXNP��*@�5�>Ez{y���@w���{�vi�z��)��2�oQ;ڧ�]pE��Ț�8$}���7�J���64�]��|dh��z���݋�״k���t�>N;R��q��*3K�N(#f�1Pbd*��b�s��\�7�0�� �,U�κ����[<�a�k�w�M���Ec�ó�;uB����!c[v�kv,Z�j;s�V�(��W���o`��;�
>q}:Ͷ�
��n�~���|��K����l �����x����X���Ϩ����L~�\��Q��T��nxf_��ɾ ���9T���ac��Iz�y�~��Z
޵����z���Ϫ�IcX�i�4�҇|�E��¹p[�S��R�b�;��#�*�pF8!c��N��d�%���n*BH�;N=�I�[�g�ͺ���`v¤Z�Ig2c�O��ZB��h}��x=&&�j V=,�X����F��}q}-��>�ey����[:0�#@'�M7J��!�X�&ኈV�j�ָ�-͑�=��"��� LWz ���,�Š論|�96>����qMqP�a��
}{A��R$^�ws�q��d���@%��K�^�d���7/Xf��`�{�@�W�m��aRm��Lϛ:`{ǲ�~ڮJ�KJ�h+����2P��l�O��kO+�<���v=�G���lt��k�ZT7'|ل8�$_�o5N�\�tCy�]�1f�723�Z4�̫Tண��-C�G��7#c��tJ�O�$:����,��M������\Gm��I+�>����X͞V>sV%n!�d_{էp�8��.�j��T�G2���=���H)K ��2ub=�S�O�_�-J�EA_B��/��0�\>�Ƥ'tCx�=DA���
x>T�A\�d���\��QB�D�NI6�H ���p�\���m{>�F;w�;y�0չ�]i�u+�k���WĪ,�!��ka�֠�e�h���d+l=7m�K;�Dm6s�i�>��o�#�E�5�&*�jy.�Q��ڗ>͆SG%�0��޶|�o���xC��Y��|f���b~�AUQc�1�A����{���Ŏ+���p��)L�!�Unx�JS1Rc�==������o�熄P,*E~$���u#R���7�^��ԭS!���y�]���d3�ߒ���~2g�N����D8�|��l�G���BX�+,p�����\�߃{l��f�[�Ǹw8fO�����f��@X03ނ"O�Fa�vnݻ������s�c7��z��B[�cZ�Lb�1�´��u~�Ϗ��I(O�5��7�P�� #<��A.G��)ż��H���g�6�*��Uu�J�r��T��M�ȇ��}y�@�ץ6��Ͼϥ��)H��[l��a�l3���Jo~�p������jw��h��F2w���urn��g&�#� '��v�b�W�^�[�g��������$�V�G_�(�p�¨VʙՃ0�n߄=Y���cR��.f� �n��7KXb���;_�W��%�&}����T.���/v�ưϥ�K��FR��Z�@�^l��o��,��u����u	�ɷ<�:�B7����ѳ|b�� K-%V�J�`���.��u�v{z̓�v��s�b� k\���gWB�=�U�8���88TX�R,bE�T�sF����S��&$7|/�^���C���#�f��,������~
�`ݵ��V�mo��d��37��f����bN����c��}}� ���b	y��!n{���>T��rV촵���G�Z�s[��=�s*�y�f}��(�\aMz�Ҝ��_u��'q���ߖ��u4�H(�"�"�<���;�����M� �6N�?TLf��Y�-�#,�藲��X��g1��G��>��,�����wӊ����%-�P%f�,c�����Ϙ��s���=r��}�� y!�[��	v�`eܟ�,�A�w
b2�؊���g�D�����m���zk�I4R�9���{�ӹ��G�����7�M�q~a�9��]Ũz��s�'�p������ �Ӳ-��ǔ�x4�%y�\�w���Ya��^g�Y�7QW;X&����w��(�7x�ps�������n��d�~�`�F��RBh-1��ц�C���C�2�{�jĐ��w���;���g�����Q��
W}���Bs6]��Ù�;�0���BD~fg,3��Q~մ��w��h�Xgk����ѭ=����f�"�7�TC�s0���[$�Ҽ��[�F�s���y�s#��ũ`K�y��{ݺ<��ެcӼ�M[���rU�`��t-�wS&�p�����+ܑó�TG��q{}�Ԡ�	��)��=Zw����C|4�G��.�Ī�}����*�wv�x��T�7���bV,���#	ʴ�G9��?��t+H�tD|(i~�Z��h�X��nN�c��9Z�&�,�#fU��n�ޑ��r{�U$]�G�W)�?p8�^VT����а,W}�LT�����_�G�Y�S�nV���6��Fuq[��^rbhC��u�s�����UrՏ�>�S������C����^���G+Vu�Z 4)EH��L����h'����1�#V��As㯀�!�0��"({�◞l�𭘏69-��h(�1ߥ�����(V̚�Am1�����R�!����U[YT*��V�0Ƿu�w�Mgm}���rRQ�+��-Pn�k�Ϭ97+j�mͮt��-93�m��z�W\9��q0�;U�\����OxEX���|7��Y�Ba�k�k$e��h�{�u#��[����F��~J�}�q,��z�}1�O,�I��x0H�'�{ܰ$�Ώ����o�ns*l��9]e�Zc�ןH��6�r���Tql$�@�qg9�U�~�f�E����l�U�P�D�[>�7��&�]d�};��Edi����nm�?E��b2?}��幼Τ�^{��,*]�鶴�3�5~�Rҝ��7ӑ�+Sʘ��7�T��5�9���6�r�����oJ�h�5c}"��mݷ�<��<.Y�y�����_�&���~!Ͳ{���)O�QbǮk�hm@�gT�5��%F��l�Ҵ�*����bBk/���n�z�+�<�w҃�u�}g�D��=-�D ��g��c��6ޤ�T����diNKm�>��%��h�[7��9�=���N�3�c��f�SE�^H�w���-窂��	x�r��rbz:��n���H��2k_GGI�OlJzxm�NOYE)|�����Wv�8��S���W���$��D�r��"���	P�R�|���i�i�^W���(�65W����I�1{����;�1��Fk�d1ir� /W<�j��r\�̓��z�5�3�h���q�<�����Gw��z�>��8�bAS-���ǇT��C<�gO�3��L��,���G;]��N�=�d^z+8Ӯ���{�߮;�rӌ ��VY(Րp@��3��yEC���H����bO�86ӈkR�%�J���,GD���\���T��0F9�1Mj�������iw?mj*ZI���(�Q6�İ�=
R�|�l�xCi�7��V����E��{�_��u����}v�����IF���!�s3�S~��/�f9��g�k)��Mrכ1M�%��7��XF"~1��V��p�C����u�����9,�<�re�߷&���Ŋ>0Ͻ;������;fL���bgq�J��|�etꢢ�v����h�� ])���,u8��{�Υ\�'�N_�l6L�[| ��;��cđJ���	�7!a`�x&�~�^��ء��+�w�f�V�i���A�~�g�v�a�6���;��m���zA�b��GD�k{2� ����a�R������) ����d�A�ĸ���9}܏��T���e%���(�S�U�#��dtC�������k��t����7݁o7�f��lZY��^�;m�]i�֍މ�*^R��Xq�A	?
��S�׭�q�T�UXْn�����oUn����P�����<�y&�Fz*�jP0>(W*hݲ�`�����l�Di��;� �&2��6�Uˢ.sv�T�4�v�L�����L!��{x4�m)˖{� ��w�	��؈>P�G��:d��Ȋ֬�iL�qm��6� tp����_vѻ�j誥�8rTm�̼���I�rˈw���*C6��0t���������?f����{���{��������j�nŝ��eP%CɁT�B�Q�0�A��)wF�����C�:&q7k��b1X������k�/0q�Z�bv6^���cw"�ٶěs�U&��C�nه�v�̝�z�ta�a�"j�,9�WB/�^�O[�p�lf��` �Ű����gX�+ķN�'�[��u�����8��j�J��ǆ�^k=��/�y��$��Nsn|԰+��ܨI[z��Aԇ��/Gb��9y���iٶ��ݷ�Z��'m[��4J��'�'k���c���e����l�P���l�[UΣvm�#���C��W�wT
E��_��}���2??�j�9�k5ޣW~��=�&`��v���Ӣ3r��u�[o��VM�����?y�� ��^NÇH7�\{:t=���}3)���:�v��f<��r�O={�m�]��_(�x�w֤��u��F�
v�@Pe&����v�Ԙ`|�g����{40����}��9sj ��)��s��7޹�b}��{<�`o��.���K��=&�7�Q�qˣ�m���[Ș�=8�sݞN����J6�n*GZt��B�6B�U[K���"�f��@%�h+VJT;W�5I�����>�uװ�%�!Sm �IX��}�V��IV�t�3��MS;-�������m}���^�2�D�{"�5�y�g�=os���S��6J48)T������Tߕh1����j��{Έ@�}9ۉ{[�=�+\�ݓ��o��}����सg�G���h,�W%�f2��#;��bpk 3u�i_�[���I,�����f9����\X��%�:5]�9����������@���l��*}/(+��hB�,4��O�Q���P�Vn�Tyn�mvwm���sZ����;r�B�N��'��8�K����k+"$����[��D��^$�Q����7��� Y�`xeG������5T���w�e�6x�-��3�uy���,ǋ|�l�Ɖ��^t�;n�W����	 #��ӘlD�!6�61. C'�Ҵ�&�QS������n��#��C��"'�7~�0������'���\?C��q��	x��؁}�e	Y��Sg9�#:��Q�|*b%�*õ��c�RS�u,��z\��N�ML򻝟�]v��F�I�sկMnc����M��N=�&�=�G=�m��wG&��sV��&��M������wv<�Z7TB�9j�aw@���_CA;:<$��55��AR=oM�c�h|�G�]�1|�2``��ljLy�]��0q.J�b�#�k>MrE�&��ka$+a ���n֥b�]fE��>��C�ɇ�L4o���ʈwx�2!<����-��K�$~�
_	8;wc|>�Z��L�DE����=��P�|yYz��W��f4<v��ӄW�E�^"�7Z�
�Ah�I#��ax lj]�5�(�^y���o��l��^�0�YT����b<NL��2D�")*� ���y5�����s�b�o�h�ܗ����jZ*��X̞�=���<��/�����[��t��Rv�K�#p���&Q�K�$߂��Ȁ�Թ�28�\��lH���n|~���2�����&�Ʃ�ȯf�5��6x@Q@��j�g5��w���s3���Lm�證�Td��ݮA�$#D#��G�h^�q�ߛ�|~S�[|�e��F�a�!�7�{��b&�|��鸁�t���S���Gٓ������_вc�Fחf�������;�W�n��$��
�h�D$Q��/M��y���ጎ���nۛ���ۤk��̝�&�v���հkZ�h����p�RWG	]�V�W;ToK��w ��GWI���
ϛC��fp'�O���K�i��2�㴊�YG4���y�kz�x�Z�pnۆ�$���S�����񏍾/��a��SY�N�A��u���)]Q��+H?!��˜��[�M���v�ɦ�w�z��|�>>�ڀ�x�6�U����0����ϛ�DW%�j�:�������N��('���1'K����񓞏J�٬��@�w"�պ�	W�2&�}zd]��&,�zȽv����jY�������~���azZOR���5�>=_�M�}B�|߁�\T� ��iO(�uz)�<W)�v���w(I������0i�{�w���k` ;,[�{�����I��^쥝�Dκ�V앂�o%�\��{UL�1yp��m���+�dh�<u���}����=T<.�GI5=�C�O����(U��7D�HM���J[�)|:fw;�T5�jv�fJB#t\�ڏ-�-Q�k�jS��j��z���h���њV�bRf�f���n�W2�GS{ڰ��H�� ��XM��v1a	j�ګ��n���x�BF��+�����On�.���O�x꽷��|}x/i[�⫧��L������>�4�{[#���]�2wZ�����h��BN���Q'`5'alL�47mPɯ�7^��;UcPf��2�����)#Ў��矃18G��3F>�C=4ݡPU�P%M�D��Y}qq���Y�>Nת@�{͊�����b2�
�9�[:���]}7�qn��O7	�V�u�u�&ҩ��o�����'���q��}�7��j�����\�F��<y��\�lɨ���[�x:�st����wD�|��T�K�Ҧ�Kuv%Mk����;�Y{C)�O���2ڦ�qt�����D���+�^���YrVT��3�L�q��ﵒi����zjº��ӗ(zE+���c�Jk^���z�=��ڧ�[�k�U�ۓ�J�&��p9��#�����c7)�� ݉U�Ģc!m,U9BU��1j3�S�UEj�R��U���<����ɦJ�ad�T�{�i������fk(�{t�nZ���T��[T��/&��Ǿ�k�4"�0�1���Cn+iF�����ּv`�Dk"<�3L�u��d��&'@�mP�1���tfh�v��Y�����0�1�����^1�.��/KX�(�%A��NBQ^V�Q�Q��.���2��ELRt���yI��Xx�1�!��c��n��k��}�*oy�76$x:��*jw�i���/�14�g�i��8�0�1��̸�q�ϵd�VJ��_gݽd�Yj�9���J5�"T��0�l�jFx&��g���n�s���e�|
c1�8�d��d���O���st-:����{߃����O/f2{���Ɍ�,���{~�p���<i�N��M2V}��SL95�<o����m/0���q�؏8n�)�ϥ���Kn=�#�<s~��Y{��&3)�]}nq��Jk�D���4S+�(2��q[J5��=7uẌ�Fo�D�"�K޺���1��5��]}�$NJ�e��
2�E[r��ܙF��)�if�4�W�$�l�q�3l����fl�6���ɧ�$�u�Ɍ���a�c5��4���UQV�ҍoWI[Q��؝0��M.sY4�Y�c�5&� ��3q1���|��7F/\�r�P����O{�Ho{{�5���
c
�1���Y�I�Fc�ĴF���q���Q�֩+h�Di-�<��e��\Q�,�+	X�3Fg�Z�g,���ʁĩ�vx�W��(׽am�E0<��nDd�:s#~���#�ž]Yߴ����N;�g`�R���މS0>*����tc�m[GNi��s$K-Fi�5M(�ig�׷���=�{S���ɸJ����H�u\x#d`K�A��u�;u�I�N��;t�..��7Y�_6z����NP��B��R��֮��h��"��}�p{�z��$P
RvҸ(߳���ٜu��>�
�#��Wmw�J�Q����7b3,6�?|��:�ww��B���y'��P�1L�~�F��\ԏ��-���ڝ��#�Cs��Ƭ�yr�ȏ��hC-�+��#d���z�m�OOo�葕4���/a�I��V�1NmM�}����uu��S����M�|e�>]v�v�y����پ�+iF�Di��a��L<M3:�̦jm�@�ν�I�Vv���3�ߛɶJ��M��6ʜa��v'L�'�5��7�J�Fcm1������,�Yd���������p\Ja�������eV�mm��+vT֮Ɍ��f0�1����}�َu��J~�|	G��K�����>u[��k�8��M�h�"K���+�M���;B�z�Xv�ɛ�!��;�a}��{�^�H���-�+ŝ��8��U�8��:��X���gz�+ia�����-q�ߋ�-v.���B�7b`{�{�!�,�v�x
��fS�����ꋈ�E4�qS�D\��I��<r9��x��VR�]�A�rje;@H?��}��
��浗pY;e@߰�b�b���Z������e�Zh��Lִ<�$>� � VZx����9}�u���`A
�l#K�����#(h��wS��Me�Ҙ���Y�wc7��M2�VV׷�2��8Έ���&�R�SH9�X,�o��&��{�'L�pbW�u�j�˥m(�ٝ�3�~.��jп��ywP��dyu�wļ�����3gr�২D�ɌJH�*18����O��N�Ns��/�Ë��3��;CCĀ7x����6>x��@v����T���5��9ݡ[��K�N^SH��M.�3���?S�
f~~[� ~7�~����ߤ�w��Q��:o�4,k�U8�ȉ�6"�"Mȁ5$�R��P�;��sF�zw=��V��=aVV����?z]�T߷"������<�&HTb4��7I�D[w�x ��k�o���̮��fx΋ap�;��ܗ]=��E�H[v�\����3qn��6�����<���k���g�ݑHN2��)m����tj5s�n�\n��N��o�Ӑ��<�y��>��.�;��Si��liu�lц����������W^L�.sۭ��P[��q��㶮�`��_OOL��س6[zF�+n �����@N3��e&�x�޶����g������o�ݴ�^c��m�+F:U�n�-�۱v���AƵ�n�6ٻWFXc4���5��um�hcvuӭ���"N'��ۗp����LBj�~ͻYB��V�o�����MV��1�չ;]�W9ho|8���轪�1���Q���.T�<��(N��	�(��/Y��b�@��<;��}���v��PS�qGž&t�t-�+�z;����&A.G��r�yVM�i�k3o�>�<V���n��M��Q�2p�ݚ
��>>�8\щ"}�B`�y���r���Y!
��Oc�7T��Wo��68�-!#�e�E#��=��k����Qr�R8�ܡ���1zX��q\���W=#�ֺ����;���δSp���Gi<p��KmG��$)���C���J���%mFk���A��j)�ioqS�A�х�Vż�Ղ�`�T�Xrⶔk�E>!�iF�F�.��ҝc���8C���F��FFb��g9������*� �VA�U$��ku�@�_j ]M{̬���ԳLH�O9����bn,�n� ޞ�.>�$��3�&���wa�I�ރ��߇�Z�H�j�81z�-�!W��U4���
���Ld�c7ް�������a�=|��$ �a4L�<���jXۀX9��ׄ�`�����7�X�k�4����
��*n�O�j���)��&?
��e�E*��v�GF��A��+V�׷���؂«*E��+�Or���R��<��ωa{���;f$5ʤN3�ьvx��ц�506�Cgs ���!eg�=rU�QM�-���)�r�B�9Ih]�u!��"k����i&��u�M�`M,��V��@Y��ZQ���F700�����x2ťƠz���3�}��F����vZIRf��3�T�M�.}�c� )+U$X3��	��z*��u�q'y�!cP���e���*7jv�[ ,NK<af�]�m4��\=����,�-�h6йp�0�#=��hx��b�b��+�Amw^4U��4sp�n �k��^�ުX,�$lC/PZ�t	��9߅O.V	��]h���䅢�ј�|������i�� ��.��91�n:���Q�q�V��dcFWou�v�K
R�����,c�xCI0I%����Cq�UN��mk1wV���,b!m�D���w�Ꜵ��ݤu�\X���}m���KI��
b4н��i��,��+�XJ�@_���ffQ;�L]�u�ق��8���dėb�u��t\��璘q��]nW��.n�:��R�5��C5�-�F�N���yX�-Q�y�̗a�a���`���X��X*��>OZ[Cj΢Z��q���l�+ ��8�a�� �@V��z:ݗ	
�-sEi�.��9��}BsV=��S�Rm-�.�>��ZX������OV}�?�Ov�b��Ey�����*7.�:��kǣ�����
��!R�&���^({A�������[��r�N��O*��4X�EQS���{�ݙ�W��u�Q��-�����m���5�g�t�����6X�,��,�R̭���볮�9�$HF�"���֟.Ǝ%sy^x\ϴ�+F�J�R�N7ST%m�sO��1䥾<�~���4F���K䬆��Sn�5q�v�̶<�H����9�\���}W|U������E�2�g鯐�s@`و&\�����+�OO͟i��lp��@�Gdz(���J1���c�;C�hh��g�w{߳�=��{����|�|{�*��d�6�s72����;��G���~i�P&6}�n[��!�+ud,�6�&`�G௃�{�=�hQ�H8\��q�@qY�>�ݘ���&b��fWG&�YB�n4���G+�����l���|�XV���E�AI��9�{�}���^�E����tG��G�|p|2�"y>j�^�}��B�!j�2��!+!Wi�ϥ_���A�mv@G����[6,����"��㒏z�!�K���/��-�x~Kwn���孕CU�/�v��H�	��5Pm���D�c���.>�-:,�n=Sk�VB���>@L]ɻ��>=����E�&_nz�r	�g����8ώW�(�b����E�����qR���m����,e��O+�csü�}���8&�.
�,�B/1tc=0��wO|{�)��͇%�z�k����`��`{R��D݌ݩ���E5Nѕ�'�({98��5]㜜�Oa,����-��t�S����׹al"9c��~�ȧ�\�������p�M�Ǒ�f;��d^�P`B{,C4�zr��;��f�%�<�:;��%W�:�N�ߗ��!���o=���^b�x��F<}�V��N��	�p�_s8fyG���A���N�X����s�/��8�.�"1#��{V�ҝ�m�j���8���/�Y��vJPWX�i���;�Ȯ�xw�;J �ͰˈR��Y�l�b��[f-gZ������b�2�%��/q�>#�� �����;�~�{���I�j���� [* 1*���`�g��Ǫ~��<Ő�ܶ,��&G�]�py�K��,�#�&���_F�O���o��m�ީ���ˉ�q7����pL�6��[h���v�[��gTu'=�x�|d�d|��#�N�L�}q�P;z������ΫWFcsZ;&��AAh�P���&������ZΛ��Z���LA\9��ܠ��V�l����U�d�c�k�A������xה�?E}�v~֤������B�G%������!��K
ݬ�X��>�ӯ���gD�����c��_ш5���-}��(��rk<Z�xs/7�XIy���y���a��xu�pg�B�	�׽�˚���� iý�y�XYft�\�Y��.�u���B*6��Ej5��+V|�$��R�a�ZxXhA����'o�n�I�YU�j��-7Ot4������ �^�+���K ����5.APQ�����|�q���ߟ�_���v�QH�X��)G�:(n}�]}�AS�o�P��@X���RD4�����f�� ͏���nT{�}Ρ�D��ԯ]�i#�UB�X�(����s3�V��SA��p��/g~��u�W,+ Z�e�Wj�U�s�|�O$���ؠ{��'�WK[n:Ӊw���W�iGܜR��}�ޠˉ�w;lI�\�6��2+��r\r<�+wb�໚�p��=�zx:���m٠��*��A����v{]FV\����_]u� �3�獧���#�[B7$T�p�ߞ0X�C����-����5����,�~��� ���"����r���::�U_�t�!��^�z~��X"8������q9�DD8+�%���s��y���WUzSew��%bcN����j�y�W}s<þ��S�c�VT�%b�j	�~c���%�ʕ����/O�*-3 )F��;itdq�?ȳ��0��*�b��څL���燐0a$37G�34s�M%��T��(g��Dog�,4	�������V�/���,��q��E�����k�_�)��te/@쪛���>L�7��.ϔ���<IJ0��2�*���*X�Ůу��R�U�@(p��.�]}u����\����ְPM��0�9���D��Ӣ�a׽9�H�U��e`�kk�<��r�����g�ה�m�I%�2�Yi$����q	����w�:��qt��!��)����VRjS���!)����C�H���	B��w��h�޸�bbOJ�og�)��܇-��y��)����W]^>������0{ɭf������;U�aߎu���k��&��X��}3�<}���S/r6ޒ��hV���Llhchf��3�X��0|���̔��'�_y,>zwI���8U�lh?B���O�j��we��Bf�Ʒ-�N��A5Y�6̐�E r�*Q��ԭ�x�v�q5��;	5��þy��~{Vpب\�9�gGk��uoNw�5�*r�ն�ڜ�eDy�ڸ쉻VۃD�g��vܥ\���;���/l���v�#k��Ά�Z�3�ݓ�vsǵ���xRpx�!��<q�Cs�%���Î���E9Q����5R�U オ�#�3cn#�Fܿ���q� ��Q�m�`w<g��ȗ>�gr��;���m������j�뷠�j��\��}P�c��$�^��J�=��]�+�v�ڎܚ�ۢw2&������4+�8�F�HI#TV�Q����NKr������tl�[ڻW��1�7��'��c��Xd���挩w�b�;�Ƨ�8�K�_�_���M˜��r���� �����G1dާ(�j����>>_i: n��oald�M�֒l)�N0�ĝ����7�4�*��!�\�NU�|��8VD 4�C��\z��4z'�����ؼ2o���pb��g,�g�ku��( �{=B�8mv���s�}�p�>`	�(�r�@M-�n�9s�.pB������y�m���+{i�=��ޛ([U����У#�]Ox���w?���{�K�,̮�epU�ZZ�����Y�1��ܳ��T�Cg��\���m�VJ�U�f�"���C��7ן}0�J���T5ZK��r˞-�o�[��J���[�y�8�ŞH��^�&��k&�M��p��z��$}��Oē�*M����QӲ<i���c��W��V��t���箭�t�����<\w�]Q�)H���:���"��Iٳ<��V|�zO��k�����Y�'zr��M�����]�'ւ�XֱVx��8�^������P�Ӟn ��!�4c���ݶ5p@�Q3x��8��^v�xƑ���L�>V^���z!%Z��%�*G�3�Տ�I�h����j4�q�\}d���:�!�Dml/��R�b�Ag�u��s���3��M�<��_�ѵ���C*�^��.;�fc��k����*>k;�h��@|h�R��� %��"���G���dO/��۽�q��U<Ω}�"j3_5ݢ�[�gF>H2G�[lnb�\M9�;>3�=��M�m;����Ѷ������;5�ۮz�z�R���뱸�_������L�!=4�֓�ae$"*�e$�����g�)��m�:��I��Z�r�N�d��bt���z$o�կK5۶H�M�ɍ�g�k��l���8@n<Q��k5ׁ��vv���&��ϸ��fv��B8 uV���3�����X���v����9����/�v�ˆ;h����6�D}i����V�Ϗ0�T�z�Æ�b������m��ӯ]�.ůisn:��r���)��5�B{�ȫ+MP�Z'�wp����fM�jA  PA�D�0y���ы��A��lq�k�i,��kK����G,����uZIm���Z�s�,S�+���Z1�٬�<�!�]�?,��ĝ"z��J���{i���Ӯ�>�^m�TUo_#3���N���g��fM���
Bp�7�H�2i��*V�����L��" D:̻���¾iH��[z�1M=LSZ�4�|o��F\?�#�WM�e����V~�M����z�h@E���+n����8�3����,m�`��m�K���I���vfv��M;H!�N:Ѫ��#VS����o-$��i��s�-����m��fd1e?wqrtZ�7���rQ�;kl�p�׹�%��h��Ld9�,�&L\,ɝ��Aӂ�	�9��K�[�wv��9�R����2��9ױ��-��s�V2rK�����x�,|6��'�|�u܅���4:�<�:"�"γ��Gկ�J>�g>7i�__�P¥x��|�^�����
��&��������ul��KS*�����Z��!gv-VE	yћ8d���&����l����ޑ��W��>��=�?O[��pf����$n1t˄W�m���y9���R�}�*�t;�7�_n1��7`��� �=Iu�?.����*��ڸp+���u�#��~�Y�3=�3�n��X�T�Y=�dnFF*QWY*{.�9鎢�K�"��2r �u/����TNn���I��Ef��6��%=��7��U��߽a�\��y�[ݗ��n׏W���\��}�[�0�`���KM�D�ອ��cyf?�fb%��a�u�Ge������������h蝥��?B�����^����g\�s��7����#&=�K��P_?s�l�w:��j��w`�^3Ǚ�f�YW�Ck*Ő`��ސ+=���}�{��A����8��E�\ܵ��V�º2�c�;{v��ݫ���Lu՞Գ���qh��gL�i�HX`����r/Z�@�REγ�p�b�s�e���ЧVy�����zb�Be��UGS��R!UF�p)m�-X4���:�Հ=�xBm�0D���HNo;�������i��]$Fu�jnhG}�0w���e���HKާ^��Ԩ�����pK;�CҺ��!Sr��"7�#��6�*�����ci�s�Eψ�a�/Ҕ_ܥ�{�������)��5\6r ��^2&��
��݀�,��.��p��	ÈɆ�p����}�X��3������l���֌)-�q��i,�a�0m&��Ӳ���ɵz�v����}#����;�{�r�;�ƼB���bi!f^9�T�;��,��1�evv��Y�S9�ȯ�OP{!��NɀY
!�5<��	�]�W����*�,K�8��D���#EMM�tw�#�j
�U��pӴ���{��w~X?e��t�&���#�T����Y�O�r㻾�G�M�
Us�;u�lqM
Z�����߁g���&|��Jf�}jC������;�9oP�9��)��у+b2����'�~~G��d�Wf�DU�%r�~��n���ƅڸ�}�蝅Bt��U�8
f���-�<���7i��$g'j~>�j��+�y���C�bi!_{�b`Ň]��0(Ed�ПB�n�/2j��<�|�9u�5�"�{JDUH�d
7����<G���P>3#z
�S�*�-q��2�VR��@�6�x�~!��[�g�`��:���w��$���3GBs��%q�.	��ۋC�{ٓ}��*!�}]%0w9��]3�N��Up�ܶ�Bd���pT7��)=��Fݠ턏\�F�3�b�p�NU;]]�p��]�7F��s���s�ӈinw>V
v�6
EQH,�s���8�D+#�
֤,����{=�kTL�����8�7Z�1�wu��~��'�y*���D��6�}���#tT���p�̺�5�"*��:���8J�`��|�3��u~qO�b�Ly��z�װ�י��&��?"#��EV,X*���_7{�&ϵ���jq�P�Û�7ت+�[����#�U�I;��4k��vt��\9
9m�ʜm��Z_������h���a�����gxD�x��]��.��ɧq��xs|�7�o�k�,Tzj�
w��"o;���#�_������>ɜp�b6�ach���rX�EF���?N�6��whx� q��M���B�]o[�d�����.���r�c�{�<�gT*�����gzr��b��1��$��[�}�NS�,-����+MX�/Ϩ^�Eke���U*�c�w=f��v�Ud�ni����-���H�/��C�O�ƔD�*,�1�;�}�y|��^�����~/�D�EUUSHH@�@�$ A��X��0�W���X�F�?s%��� � )�"�@R@$� 	c ��$�R !)O��� a!I���sBI�)	P��$���7�"�R ��D�AX")δ�i$!"�M��� �T��,1dDX��Q�*�A�$��EBI$R�d "B#!(
B�d$bIHR E�"�Y	 � I	Y$� E$��I`���  ,�J��+$�, Y"	��
 ##�!0I
� "c$R)ie<�(�j$*H�`�R~�g����?!G�+!!��?�����k?럧��_�����2�fY�����^[(_Ä/�8����vgi	}��֗>�����?$�6������I����M~g�_��#�"j9H�O��@�~߳��_���?�BB!S>?���}I�Bi/�/����A|�/������ �c��~��} ��L��������IkB
P�E$�R ��E�IHH��� �H
HA@�0 ��@ ���D�BB(HH�"�$�!I$FH ,�"�� "0�,�d � �� � �H��E�XEF)����P���$$2@��I ���B@H0�)d����H)$� ��$��a���)C�I��/�O����]��!!@0�ҟ��?/��g�����	���}��6(/��>b� F���@��_���~��BB��`P��������ܾlj���'�~?�B2e%�?�������`?�m�~���b����>�	t#��%�����}���s����� Ⱦȃ��t~ �����&�_���>�l?`. ~�����[b_XP}$BH@�������� ����䬱P�4j����K2�}Ơ��n�d�	:b��~����H@��/�_����>��Gɣ����.��TMq?��K��P_a�>����5���b���A����$$ @�!@����~��BBPa #�.h��ؿ~�
��lI���HT�|���}�?,���F?��|(�5�hBB��[g���a�T�L�kg��	-0@��_J���_����~�CH@��
����ԀF~�yHH@��}
� Q���D�k�f%_��3��?S��1w/���"�(HX� 