BZh91AY&SY�r| �߀Py����������`z��vp �Xƍ�!��zhh=@F@�SC@i��(�2d`120 2d�b`ɂd ф``jf����)��� =M q�&LF& L�&@F � �$ 4*~�)�jji�OPѠ�h6���$�`�i"F	!�Ob�It��<>�?�!���$JC����I$Ш���ʤ����]�%~�x	<n.��Ƀr����o�;/��.�=U�nz1�l;Y��U[\-KT���0#St%��qZ�&UqCnh���[�3R���i�O��U\��Xp�<,G,5[:2��/Р�g�8���VCʓTXn�ʺ9ٜ���L:�dW�qDD4	q�s�K�l��K��<���Dx�ǉ�H�j(�"=(�*Нi�M����(�[&=#5�3�S�u�f����ے�eU�UWM9�%[���s҆�S.%]��.�/�
�J�3Ty^�e{�N��5��I�W���aa���)������W��"a�+�P#W�۱t�0�����⃦�S-�b$�&����@PQM(x	 ";�0�����U��W4� 1�P<�A�l���[T2�_Ue.����&����H�V�nuj���#V�A7�C{] ͆CZ&�c�敨$9."�sE�HS7���v�1t(r�9����j�U/m��T�,Х�l3*��'p��(K��M\��%`	"�C.78�v
`�b^��9����T1�K9*��F�FoJ��buFkum�ڹY}��y���\K�[��3��թC�]�gFՊp:��v'��_�7b�k���a�"�ԚX��.Ճ�#^�$̈n�+���6 ��UC�C	�V] J�R�iHhYS���v3,��J�:���x]]��|�W{�p*�p��� "*.�ҍ�4�݄ti��L �Q���Ϭ��TB�Y�3R���^'6�f��h�{}_W��R���%UA�%>$��
��!N��y@Iw�2�k
�
K)Ԓ��m���*�AAQ��&��7��S�E��e�l�hJJa�Oq5�
%����ݜz�Đ"ȳ�?��K��hQ���7xw�� ����������"K��a�~�U;$�p�7m�.��X�Ra��b$�Sw��f���}r{��O,$�	=�4X�F�E<����n+|Z=�^�&�'���o)'��bk�o5o�*i6�$)�5Y�B���[U�u%PFa�'����ý+����p�z���+H������%Sf��������P3�j&�c�C���u�?�$ڤ�	(�{c�ka�-���)+�m�,��q|��$�T��=��E�]�KNr�g>c�ݶ�|�%ɫ&I�����qt�?�U�XW����ʩ�K��/e?��\/��˗�s)=檉$��$�q|"����Z�����A�I�b��M���ZГFJM�/�$��b��#�|`\�3YcD$�V��z��E3��l��$��.����k9�%p�p���viMr$�]c��z�==T�h����ﱋ�C�䧠ꨛ�z�>6ihI�<
Q����y��6g��u�S��©YҎ<V��r3�˩M��[-��&aH�L��!���$�cSG�j��*�wY��tr��m��#-$�L.mX�+G}��ƶ1JD��Ǿc��C`���dg��b�	5���8:��d��қS���߁�T����w$S�	 ��'�