BZh91AY&SY@ӻ�Ȋ_�pp���c� ����b)>��     @@                       P
  P   �                                      {�@( R� UPQP*J�@(
�����
 �B�P IB�  P@�)@ .�       {�AE��V��g5����h���7����������� ��н�ݛ�9�������q���w����� w��e͡특a�T�	�̢���^|�/��c�cp �e�R�c3���J|mJ��9OR���r�ԥ)����)BVYx{�H^MS��A���|M()��AT���       X�� )��=�)JYi�IOI�yt��)C��;��h�_ ;<�*U�^�|y�J�3K�O��*|�U{������<. =���dc�\J�f����*
��($
QZ;�о-R������)O��ޥR��x��U/-J���zS�iU�����T<8 y�yT)��>��O�#����/��>>�>>5��HPW�      � �H����U&��:U^Z��[�iO��U����ҩKﷀ����Yi��u*^FOX���C��y�ҴՇ #�J�17��{�)|�W����UJv�<=_-JU����|A�> <F�f�q�mW����`��[�ƒ w�w��X8�t�0��^M@�8�T}I
ID�       �*�����p ��>>�f��j\�Q�[�ͪ�����ܪ��}��_3#�k�)�w�� NuRͣ޻�y�_%AJ��Q*֛j )O}����.�C��p �`�j�؇��ydQ�s�P`��*Y��r0�n,�ٹ_!J��)B�� �    �� 4Ҹ }�S}��>{t�5����P� Z��i� >��
e�WӀ��Y�}�) ��J)]
*�}��fʁ�F:,[ǻ�Š�nl�z��������$�����w���̾s��x         ���T0 �20  & Њ~�$�J�      �B��J��h`#4�ш'�JDiT� h`  '�R@��       I�2*�i���f�ɡ ��=Oj'�:H{����'����_�w�>�C�}���	$�g��I$�	H~P�I'��j��v������_�U��l�.ukQ$���?��	$���BB@�?_���߿5��X���3���~�t~�}��LI%0�<��?�H���W���{�bzwo!f�ٲ»�@*���3�����V����gd���ɽ�a9vgZ���U�����Os�{4n���l5\�.�j�ԭݫB9���W��P�)n�>���n� �6
��m]�V��#qdӜJ͑�J����sts@ gd���\[�����u�{#�Z�m̘[qg`*��Q�d�۝����cq���1l2%�㗮��$�=L��/]AMR�	=��\�G��	gw�'s�&+ݝ�����B/8z}f�Y��c�2L����Nvs��Er3ZS}��ޗ�Y��x�Ct+����cdnM��V�mqb�����"X�yHv%���:w�s�u�B%��f�E��ϜH�T�L���{��ս�v��+�a\c�^%b����.���{[̃'�ؚ�T\K���n�]t���;i�7~X$�@��ttٗ����w6<i//Gc(�a�t�#�N�D�v��.���qݮ�Y­�A��&�b�̜�d��b�QnМ$m����u��Y�����ݗ�ot��V�m�M�n�1�`�(����{��4�x.�F��Gjܳ�WmX�4�B@%�z�12�sݺ���_,�{��`.}��|9<�ƚ:�#RaP�sj�2b�6q(�n^�qw��$%Q��	��Zd��)�������nj��� �-�C��60����8��ɐ��:b�xo,���s�S��p�5�OJgqZ���I��za��5�K�՚���9��&��a�� ��w(x�w<P�L!��w�xl�=�$�t�}�j����{��w4�-�	$̈R$�����N���n���r�4H�r]��Mi2#Yas�@NT�'K�u� H�@W�ٴ+��el�7�6���E��4@��Z��/A�Z܋%���Wz�Y�{v!%.���ӹgQݓ	�-j����0��ĭ�#	��ʌU����o+wq�`�����v@�J#k�z�
!u���nn��T'�T�3�L��툩�tT=�3x�u�8��P��#8c$Ve"XD�LQ(�@��e`Z���Z�Y�dќ)#��0fژ�PXoey�M"a�nh�;P����n�q�hy6N�1(��c7�����F8T�{�YC(���:ޛ&[\R���Es�"ҩ;��3{篵�W[��ƾ�]F�؏n^�9�f'۳UC%������͚.G���+��y�^P΂�`��0��r��ٕ�}�B��]�{wK���J�JR[���8���1�0)��c��7��(i��y��7[�=��ꡃ�_����gC�\�sp��=ݙ��]�%"�h����0f���`���̈�L:�o#2`�ry!����a	��A���#��**��!�3Py$�R��S�tc`>J�h� ܉�Gt҇tq���˰`ZY�0w]4��dD�p�ݍ�/H���mO���9ع�����ܕ�g�$������k���#X��.!�s;,��w��lxB�޻v ��{�T͹���x;�Ub"�j��7F=�Zbk�f�Y�����S��:���sp�c����r�p��$��{�6�:�O�q����W+or�ܯu��#��	���
d��v�Ϧ����;��K��;P������!��7{9L-մr�6��wE۳�l���qS�سu�!����� _7z�t���t�	������sNi�L�E÷�K�a9>��N�_v�s��9�у/|4�sFA�Ɍh
e�=����tl�Z�˭D]�0��ׅI1�jK����z6&�]���B��A���^��#j� ����V�1!�$����k�����'[�.���,ޔ�\�Y���б]��d�6�A\��ܜw�ي��Ԡwx���m����\�4s��ŹGN1�;U�;t�L�[h}J�z������Վv����sy���<D�*�r1+n:�u+�$�M+u�g��Qn>|�I&V�ns�g!´C\\ir8v9�X9�"���fn������%ydC�14}5�ު��׻ˬs�����97	/:�8������&	-�K�A�a��G]wI��+��9cn�����x��څm��䄝d6�އ�q����.^=���0�A^]B����Z ���-eJ�2O�p����Ma���D�&=罕$��S�>��R
��k�җ�K�.�k0®k5Uٸ;�;8�r�]�t���V�dl-�sy�f�ͰIŬ�-��\�=��	�gdWL�Fװn�y�Qmm}�s�[��o�uKoi��X����b��jE߻��8R��`=����(�-�ϰw,Gj��*�;���r�:{�t�ׁ/n� ���y]`�:[��1-0J;繻.u2��(����M坴'iLr��!���Gjz�;��y��&��+ܼ��Xp,Y���M}ɰnQ���X�H�%�.�&���Jݰvϝ�����2��g�J��Q���Kو��,➷j�P�|�C��ΗK7t������yD�[7�b�d�c&�Igl��V1l,�����X���뉣:B��3�ν^��� �V%j�$yrx��9��w���6)-����Zw�l�7�۽y8�@���&�8�>������˛m͏�w�DnNu��ci<�L�U�H�%�x�c�)�vl�iٔw�+Ԥe����wJ��Za��gq�����Vo�{������n�G�9�v��Z{d�z�����#��m��\'����d�6�t`�M�0LR8��>)��r�j���(�����G�ч:���Z�˸�EJ�FӊZ�m-`8��ͽ�����[��O����j�8�6	Ѻ&s��i8Uݍ�Q;�)Mע��ʍ&�Ԛ e�2c�E���;nQI��j�k�Oe��S\㶷϶B ��Z�:�[��ݙ�S\c5U���ܣ��k+J���܀�5��;& �.�;s��"��k]P���It=U˳.�,6�ݡ���Wt�z�ܗWp�J@��vw �n��J���hh1�}��V��H�F�;��׻�Y2N����t'�1Ǳ���.zwj�uҦw@5�4�hRq�`��WAi]�B��]8�Ã\).�WLr��ָ�:����� ���,Zj�U��]�7��<�����; �6D^�u�ݒ`(�vwIv���wT�w�N�oj����w�i	��W�!��P
O'�����8����
.�zFѰ���)
Ƙ�xtnf��w
vm�1�k��|���;�`5���!�Y��ar����'n�6!��v���ww�.�sw�����"]�����Ŗbg{��z�	��n�"��N���o�[ҝS�Vlwe�����CEcgh��m�݅IN�$܂=ܚ9z;��6%a�I:�ac!D#�t�޳��yK�y��B���s8@�������}��{�)�wM�����xxj��n�����	6�!ӽ��/e�F%��m�����Yҡ7��K,��Lkf��0���$2�h�.8��n�������.ܫT#�J�E����em���%7���6�d�:B�AD���0ϸ�lri��C߹2��8�v�f�1`�2[ho�{�y����k�ف�/��u�][�g���9K�N���	���4�%�8�kF��A��Y����B�h<Z�G��5��Ŗ�h&WݻQ���ݭ�kH䖩�I߯��ϑx����ኌ�;nMqk�C���[roG�T���k�Rp�(�=����r՛Ǆ�{��gLJM��D�'s�K;uwB��v��O#�OOP��E�We�.��f<��1�A��.^���'uu�k�X�f��Wx(�vg��'�0��ta��M���[�WL�M�w����w&Κ��4�鍣�^9s�$�n�k���Ʉ��wu�AY98,i��g7���������L��.��A�i*��s�K�"���jXQe�F=d�(��	�ZR���L:��szx�%U��/k]Q�5r���r�6>�p��w_�,�\�k���j����4��a��K��%ahS��p��ъ`g4���n]�ݬ`�q�0�A%�T���Ȝ�m�fQv�m�ý��ݽ̳©q�����R�&u�ZA�Ž�GZ��i<n�����#ȳ��.vt+r�ln*�b�9��l�Iփ���4$�{8-G�)��a��r�p��vg9K�yO��$э�uqkZ7���&���F���<"�5�v`Z���2Q���2�8����s1���\�Þ&{;VU�׻�=�*U�ar��gџ�nNܪ���U��Yr4ۻ>jaޜ� fJR�7���B�˃8.	�53�;�n�9��ŋzn�ї��Wzq���i3���"���hZ�-��˔�n12��pZq��A�]��Ѳ!M�ҡD�l)��S��l�Ӭ�G��`�{l��N�����<�ӫu*@]G,#�p���������]�ڷ�J���{����D��7���:2�Cyw{�#�j�ώ���d�Y�����t�1��V��yHYu�]-i�{�Dwl�r{�5y�sX�s{�k<�v���wF���;l�s�bnEA�w}
�k���Yy��Q�ؕ����=L!%mQoS�5`�sgu��u����+��9cd�N.2�:��z�xCA�RH�d��U���6���ۓ{�ۛ���8�"�����N�`�L���b�D�m�ˀ�çnk�vU	�w�oS���7�-8�w�&o���b��\�v{=au���y��1R��m��|ts�m��h��Κ
��_���� ����nE4��0"�g5�{^��F{��~�S8qqv��0Թ�
A�]��H������Rp������ޙ|�s�MJpٽˡ����ga��c�wh˗��.�#:����7��E�`�=�~!�^�|�%Wp�Jr�7y�՚�OR�u�(s��=�H:��K�CfU���U�n�][�vq�^�oLV0����&�eKZ7����ヴ�`Gyz����篶���y��l��`G�.�S%^�ח�wG�e9�V�L��&���R%�Y� ����Fq���G-�gc����vє��n�#n�9���ܴ&̋Fm�p����v���b=��_�eWIn[��
n�_i�]sJ�7�͸ x�V������!��z��WW8�bi��CY��}��l��`��"�m�7N.�˹@ں�Zk�V������`�ׄL�)�;�a��b�N*@�g:E����<+4u{����7Z�%dE͡=�{h���C�EwH�7�ou��ER�y�<_ �#r���r��#1;��p��\���6W%�[ɵ����O�M��
s���M�DKNC�4H�EU�����-�x[�R��7�Ǽ�wt��b��8��3�0��:
�#�1O��M\�����f���G6�'m�[@)=�1��ќ�u@�dD��s5��ή��G�{������O��wd�4U1����⛽����At�m�d�p����\x�aM<Ass:,� I�<b��I�,�b���NA0�aV$�t�9p��q�(���/H�o�:e]�h݁E���wN�t��n�^��=�o
Y�e+
�m��3�;)�,H�r�{.#�V	@ƣhq��qnN'93����`غ��h:�vm������OP������Dػ�:�	�`D��<è!:�H�P���k�R�EM�m!��R�������tp9��<��&\ݝ��b�v���CN��޸�(��Q�אΙ�dڸC|8��V��%�6�0b\��Ǽ��%f�����"��k�wb[�����Gk��M�җp'�t�휗7F�zo���ׯ�7..; �L������|�q�p]���$��:�]�ν�ٺ�e�xn:z�bb�$��%���=�Pq��%��^���;0��@�F1Aqq�Ct՚�0�-�Y"MRp��,���k��ݒ,��g�[�oFP�˛Q\
�XD;E�ŗ����h��q�{\�ꈧ��9=ݗ�U�U���`�8'>Ֆ��bePp���R�x�T�կ:j�ߐ��.뺅���v�T�ƺŽ�wOf�P;��6�+�EŅ�m�t/N��F,� <�4cdS��Xl�2�jdԩ\�npV��&j:-����9-8�[,�ׅ������j���n��j'T�����`ÒF7l�����JB�y"�6�ڲ�b<(�\���O_���N�5v�۽�ގ�p�,)�T��p�q�����{�syn;Ӟ�n�/g.▘�I8FqP6L�߄���u��i���u�W\�֠�V&�\/狻wX�4�z
,r�����Z�/on�ҷ���P��7{.�7q�|���vLծ\�k��6��غ�M؝�w�K]������(cfoK�Y���3{rL8s����gܚF���ZD�v;��2�͋����Euh;���H<Zy�� w�Dټ�~b�*�%����rW��ழ�����M�NJ1^�,E����!�4]�#�ݦ��s��.�6F�s^�7�3�p�΃:aG#]��o�.���ˀ�+�E+�5Rb��Lи¦r��<⠴��([�����z��2� N��&�zIR�.¹(�ޣ�n�z�J�+Lt�H�ڇU�67��[�q�jV�q�� � ��~�{낪��׺����Z�Ɨ�K��n���~���y���{|`�t�k�u7K��T�[����U��u6��nOi�r<竵R��\���������G�����2e�6��
㳑�Gݎ5n^7<F�M픠�lv9�4�-����p�G���hz�jon��k���6�Ź���v���)sv�v.b^#A�ڱ��m�iۜm��GSj3�y�:p98�:��Z�sE�t*��z{nn�:;g:m�;�����˜pERn.�8|���㶳��[r�[qs�<�/b�g�>�h����	��gX�[qՙ����Ou�Z���s���܍v�u�6��R��&�6-��4��o;I��8N��c������ta��.UK��۲� [�k.(ajs�-�Y]�G�ѫ�n�zCer	�m::�j�b.*�6�.�v*����]�Q�ݢ{Y�lx�Y�[i��:�c����6�������z\���u=gc���F��E���x��P�z��]���a���9�S�y�v�G;hԱmASdKn�:�Ƿ^ku��2=�#v�`���;�p;�7ki�Xk#]�v���8�3�>zSv���j��2��*pk�s�j����Ƭo�G7���۰���[o�Is��y�n����g��=v]WF��՞.,P=Cv���qu�3k��nlv+`'uz�kZ�Mǰ�q3��=�ù���+��(�é󥷠W����
����̠Im�L8\Ģ�8����Χ��󝛧�j��m��3�T��t/O[Vmc�v� =�4��r<��^;z���4�{pF8ݳ웒Ƒ�Z��m�����699�V�e�8��6<ri}��ϛ��\Y}���Wc�K`h�ƌ�,��:nW���!q�T����x{�
[O��p�w&�u�x�㓆��L{:�<�s��nV�I��7)�p<:�3��̑�nvu=��y��1�KJ�\[��m��'�"��v�O4GkH)�F�¹��%ӎ;V��V�.dHꝲ�u�Vs�l:�ܛ���s�U��}�M�d|Q����6�\߇�u�9��ľ�f�>�]Q;%��T��A/)s[��Ş�pE��:f�)��\=1�;n��!�� ��u��S�m�tq���^�*pr���}�����\�r�y���W6�u�$�u�κ�0y뙶t�M(�1od�瓏eg�@[ 'h;͘��)ѭ�{>�qe[��������w:��]��F���y��۳�m�ڽ2�9���<ι����w=���򒛳c�A�b�۞�u��Cu��b����u�Ǯ�N��=�g�n�{�++g�ܼ�9����L����{9��2�vEyŬ$��똻9�q��u��9M��{���m���pv�j�˝���P��k�ˎ�XѫWd;yF�[K��[Ip��n��]�`�w>ۮ3�x��m���p���z;���z��zPS�[?ﵝ�m�4�G!2�n���ɻg����$���q�vl���b�J[B��;qN�B��v\�_p�M����q�|:��[�������I���.u]Q��nwY�8�3��"Yפp�]q�cצ^�֒C=l�{F�q˃���[GF:�ƃk����Mn�k�m�kՅ���;���I����cH�*2g<�^�[q�e{>�����8�C%������]T[�Gj��n͏p�:����ڵ�Ь���q��ͅ���S�7���)=f��n;-[wm%�m0Uۧ�Nwn�q�`�({6;������d3��¶�qӃ�\��{g\�=�1��<�rv�:���[u�wMh�ڔx��U
�5Ǡx:]�۷(��r;��;��F���U���tr�n�h���:✧sr������X2��nmۗ���g>,	�l���\�Ƶ�k���27Nђ��P�|���D�K�N��{0=�5Wn��c�v%��7�����6���vW��;O�]�\�`RU�:�b
���33u���4-; �tۍmw<p���մ��<�Zz�j�{C���.C��vz��:�c0{nN����åk�<`�0�h�����A����/$oi���=��6����#�^�8�큓]�ĝd�w5q5s��`p���h���m3r����Ƹ��ǉyN�T����B��vW��=P�r��>ˇk�v�@�����tyl��}tt���7g�r���Ҩn���H��س�2�哢x����˽��La���٧r�c��L��ό��<\=��t�����d�l�\m�[�Ã���[����I�;�c�7"��\
��v9�����*���n��Œw�>O�e�*ӕ���ؙÊ�����,�/[��Ůwn�ذ�ӭwg��<�Ѓk��+�מ�O�[u=����hq:���u�n���e�le��G�N�GV�����8������.1Ogjm�<���<?[��=]����c�|�����4r�#���E���<�c�o����SN���q�����+\r�Ṷ�/Nv��<�p=�2��6G�9�z�0 ��k�Wb�bތ��l���s����z�}^7g�jʁ��yܧA`0�W�uz�lGZ���ƻ��+s�#{=�O ޴p�f�v5������x���B�<�����n�O��I6��e�]�g�.nw%U�DtI`�v*����W������9yc���t�4z;s��뵮��q�kvP�}�í�n7/%���[T�����?8����d�ct�����iu�mz������o���Cك�f8�j�i]�6��X��7k=�ޏ���e�{ckF���{<�]U��N+��om1<�Og[	�{����s�4dN[͝�+s��q#Q�񇮫�u���3��ev���-�m�C��*!۰whxFH�cv� ��/m���9N	�k� �(ȇ�0(x������n�wo\��Ͱ��ё�nxz'��C�8{Z��[��[n�ִ4l�+��m�pM�n�s�c�9�d�Z滷]�Y;���DK�H���\��]'[T�)�Ng@1�	vh�چ�љ6�O�F�^�-�n���y�c��َ:��m��:}�,��v�.�E��dN��e.��D��"dcX[1+*k(bE���Ń�<��v��1��vN�=�ct�{e�P}����o�,�+��:��C��[�=�>~A���l�u�k���;wV[��lc�=G]�Z�@B�@gr�3���rt��ۥѧ����U<G�r�ixֶ݇�磙}��xpk��'8p�[�gm����p��A)�:k��vzG���Pv;74��vt����rX�[�T��0�f�o��K��j��u���K��cS툐��7%�:sZ�h�>�"1�J!��k��ۮ�����Mqʅ+�9H��w=��Ÿغ�l����w<g��z�m9�×�t�s��k��ˀ�E�p��!���Z��p,ٚ.�D������Vz�Z�d��c]���6{9�����e�8ܘv���(��hˠwN��*��~��nnĘ�,V�����
wFs�^<�%�1Itzz�l� ��ñ�燳s5/E�a�q���u���Mm�ר97��A&��2��SÃUα��bm�"��j�l��7\)�����]p2VV����σ�[�{l��/8wJ�Lf��d��ٟc��@on8�����l�`
K�x}��$����5���0�ě<�n�K��ۍ���ة;k4������ȵ�:������)3�Ku����XV,.���k�D~=�8����������'8ݻ=;�S��m��2��0V�ڐA��q]q�ZL�N��ۃ\=u�vN��{7}�-��=Z׵A��%ݒ�zy��/: ;���r&9�{����m��ۜ�V���l�a���S6��N���^Cŷ���Rn���3�nκ
$7�L��v�Z�猘z�s�	g��u��+[l|ո�^~��Ȓs<h�<��<v��6��,Ν�������wgA��x�ڋ��+���<󫠝qe5��]��B^�#�]��P��۟i�͎m���5G\��qs�ػF�w�MFyx�E�j�-l]�6�oh��s�>!:�wh�A�W	�+��=�rm�3�+�\uюݎX;;�X���9&t��m��&��=�[�]�m��V8..��v&Ūm���k��V{�=tkp���g�!�3hq���n#k�g��z���ы���Б�)�u�盵ڨ��8� m�fv@��s굃;h{-�I.��v��F��x�v2p�n^�C�L�m>�ͭ��$�>�r5x�x��y6ה3�:�z#=���ׇ�-۞��y���.z���;bv�n*�ߛ�v�n�4r4r(��qpi��ݱ.�$pM���7[u�#[O>wO(mcw,��|)��]����v�;mF�Rk��[u��n+�GN�nv���1#1>�űU��֥2>�����q���ݗ`���W��Z��]�[���8]q�rn�{+��<���V���z3��^�?6����b����s�jb5i�;�Eu�>ldL� ���m؝�L\�s���`�$����%g�ppv���m�y���s�q�v���kxI-��V���*�waޑ1�,�h��"a8Ͳe6�I��j:�ܧ
#�)���|o���v�r67%��z��v�fwI�v-u����-־3��C���:��G��ۜe��eU��m������'H����l�#�d����	�񃆼�]i:J٘I۠6���y��=�V�-t<F�\�4N;�v,�lp'[ck�-ڸLm��{��Յ0Qk���r�	Hc�6�u��6�{t�f��K�֊��O]ۓ��=#���I�e�1^5��-�����n�&��7G<WTh����v�x�属1s��C��͉+s>�(�����)a��ag5@v�:��۝�'��F�ɴu��	��Y�2��
��^0��..��z��'g��{���rv5w[s�ޝ/u��b������/5l�IL��m�K�wCa�mHW.�&��<[��N���ۊ;e�Ɲm���4h��&g�ى7�8涬��6�i�3t�p�nY�FΞͮ{`���k���fη>�>v�u�Ò3�^����\g]���M;q����ohC�i9.���^5Kq��n�v�;�����kU��:�iu�_|�>�Y7��囧��-�.
	H�ЪT*���($�gZ����?������~������ι·�3\�;���q���Q�d��iz�h� ��;Ś	^�\��·ke�0���;_yzt�)*�|���{Ǡ��*��l�Pl�7�2tc��1�	���Yf�o���}x�R���^�:,��:��:�C�ĳ*P.0�����j!��96�v��:(7���㐮+�NٗU�=����x��>�!]��u*�U� ����_xb��_E��˞��LKN麤�v��ܳǗ�{=�����'��vΓ���&��+�ӗ�	�F�Bٛ�e�#w/�:�j����)���Zx�V�;p�r
Ccp�^��%9yz�A<zN���S���C�l�.��%-��_^͹=�����M;�=|89��?_]�v������kv�3{��O�Ki�C(�#��[��_t������>>�U^�<9՟u�˚�A�m~gBP{y�>�L9�4�z�¼z3���&�����՗��^˼>A��H�X��e�ż���Y,�yXJ�{t��a<\Z����#�;m�Ç�l�G�y(H~��ky0+�|�S�+vCg��f�z"&�3z�oa��`���5$�����3�j��� �^Y#���k��q@$��-��]��k���¾Zj�tk<�����H�S�5�,i�8𸣧h�����;~�Vǭ�e�}2ވz�Y����S��e`.�j�'q]фdNV����.�֫��ٜ����#�e~��݃��-y�Տ�瞭�{j�>K�A!�s
5��Ԇ_���{��BWW���@��Y�VN�5J��͚(.��4�'
�Ç��>�V/<6y�=ڭ�Ka�����ޫ<V.�Y��qc�9|5�}$�tu�Og�ðv9��}%�=��M {z���M��@��}����,�����<���\�;C�J#�.�mC���r�%�������[0�S�pH�ɂE,Y����*���l��_c���z:w���D��\���[�ܚ����a'zT���(3WP_Zd�.<g{ݷ�U�qK#��g=��������3��S�5��9�LW��ܠ���{V�xZ!޾�S�*+�5�ۃ��*ǜ����uN��ϫ	���N�n��r+a�L^�q�=/Aɋ�j��]�{;�NxN�qd�WB��5�{7瀌�����N��zo]�uw��[��$��sr{9[f�����qm`0xO/���a����6��3��.�#��,�{�� eje������W��鱣Yd-�5�]#�!T�!�k6���59Y���+"�1����f�5��5ߎ���N�� ��f34<^�*D#���2��,]�]/��$;��l�O-�Ot�ə״������*1[��= �};V�D��.�ܗ�s��N���C^UF�e��]g���]��m���AѾ�X|sػ��s��{����p�B|���p�Ɲ��[Q����z>Ǧ�+W\��� $�VbQQ�4{�零���9��,����"FV��n�i��R�����{i�U�_A:�n��P�ع�xB��yxʳ�75���X	)^����ȫ�9�_�~��dxx�u�"1�tv�u�8�=�"&����Pq��3^��Xy�;Ss;��ot�VᅋaF��ú�{6}E�{�$v�(�}�(Zi⃓����F�$`�jovf���'NLZ��������}�*�)�V�-=�����XE����s��&Q<�C��T���خ7�A�F2�U�ڝ���8��L�ٽw�T7��E��x��2I��t�'8��l�Oq���i��y���ܷ�q������g.�
sP�����;:�9qS��>s5ข�۞����p�E]�2�`� �lKoF�P&(C����"#z
I��5v�^3ȭ��v5���;P��k
�S���<*��s�9k��m5���1��o�a��ٝ���Aw�����֘�&�9��:��rR��o���ټ��v[����-X��ۧz;�
���~I��w5�B�������`�6�bR�&{��I��
���l��8��n��$u]gQ`���V��tQ~m&�}E}�>	�~Т�ʐ�ONK=�"K�0�!kHl�b�ÑP�NQ�Y�I�|�s��g��x{L��]�]�"��K��^��L����H�p��;1���.>����xy�}�=�~�D���hAc�I�rY��ۦ�7�'fQ@9�2�[�Nμ��o/i���4[��|��_L�M��y�o���4�����q���+=�rz��iy�J��y�(���#&�^��rgUeFb����S���T�ޗ3�<�OӼ�٢o�|��]�q����������������e��T
<H�~�V�R=X8Ni���}�t1U��|WFr5����ۤ��I^�����nw3�Ѹ֎y�G��n�6YO_�X��z}�I�n�.)鮋�*��V�M�`���D+jŮbU��L6@����@��B���y}ΆӻE���ܫA��807L�I(cS�l3�4�'sv�H-=��]{B�j�&�P��\�'w7d��y�2N>��:C<Nxm����z槾)���g.!����=G�tP ��ͩ[�7��-����I.$Eh��9�î��'��������Q��-��0״d�Zs����3Z|��7 ��}6l�#�^�Ue�23:t `�Ҷn'V�|����|����ָB<�sS�����S�wȧonp`�-��,h��q���Tfh�P*���aN�&e��=����4���`]z��r�SîqZjɽ���y���:��z6�X3�4�oP�1�e'�k�l���U���!�J����ޯ���{}%��x��#ٓ��{{b�Zƽ�/�3��;��D��s�t9C���{���7N��}�jB#��x)�s������WI�{����o������7[�S��ܾ�=������v�M�� ��\\�;�9� ��i۳s�X=͸S=<�qo��+\�޻���5���Y-�sv��r���{ne�6ˍ&�*��ܜ�3v!f�m���R����ݶ��Ӌu����n-���V�����3�'�A�6�L��=J\���6���)?�=�=���}P|s�f�_=+�$ǻ��ά'7������Y6H�`�bb�*���F단!k)���C���|��=Y���vu�~�&ԁ��yn��I���.��8Frr]o�ʼ���u�ᐯL� lc��w��k\c�e��]ll�9�WՊR�/>.���ݎT�n������+�5z�HQ�)d����D�cHꊬ3|��z��x�$����A�+}�ϯb�`�c�g<(yg��\�vz,D\�����A�#����l.�+����#w�����;��vw���uw��BZ����>�Kt�<!�H����p��e+�[��i�+R��0w�rf��݁X�����9F���܅Y[7��B���A`ḣ*V���@&�	��������<׹J}�\~k|���ZY�#< �9��EӾ�H�K%�#�,hi�y�5��
�^��P���՞��\����\�;����ڦE��þR�7v'~�s��J�ꓝ�W2��Ѹܘ���k�Q��wj#wfl�����7c�{C�u���K�3��3��zL�Nu'Vz��{������@��J�e��E]��M�kRz3�6���)ى�J�n��t:�{:�ݣ�]'�s�r�sׇ���¯Nz��]�{�1�,Ѯ&V��6*0�3���%a�*��[`�[��)��{�a�Mۋ1��<eٙt���T2(a�w,���T�8nm�˓�f��X��3efD�҅�(�!���܌J��+(On����p�>S���0�k;�8����~�Q��1��U�o��Z����Ć_=ȑ�yv봼��Gܰwc���
U	;�0�O���I۴Lx2j���-H����p��{}s
cb�:�^�b6kp\���XV���cGc'��%�g{�+��l�`��'��7驾���cO{��(�p�x/2��Q�<����}W���b]����Z���ǎ��漏/2Ҟ�<�HX���r�)y�[�̸.�q"Z�m̛�w�h��&p�p
'�񳗯������yE���Wd�Oqz��;���r�׻��V�
8�_Y/?"�*�N� ��`�b�^z����:�K����C���^���5����d{�w��xb��w��<��^8r�&�� ��c�=��7�O�w�{��o{Y��3�^w*xo_qû�g�*�9�+�:n�a�l�Շũ��'<���ݑ$��ѹr�U;�����'�s��>�N:�����ł2��/C���o���P3�������/����EF���oe�_�m�ִBqOU�z�ef�@ܳov5 ��ɋ(M);HE,ʸ��^6Vh9j�R��=����e�>~"�1�pdM�ɩ����:�sl\��.sSx�K%R1[I�I6�uJ��!��n�ުW<2�o��Y����V��7V�LEs�7��n��{��s�d� �xbhNxYɻ��y���T�Vm��iH��pL<�Cwgr+lj��q�GQ��n�ŇED������W�z���ު����|�{��>�\��{���3����w�?r�FN����v�o�'��i����u^�'j`��X�-B:/d�����CNQ������Vm<r����&=:�{&�O�o��Z>��ΚzR���霍�Nv�����`�r�)xPޝ,�Nz�ƍ%J4��2d(�f�$���O_&���i�軙:k۾�PK�:�U��gA�f�"���2 ��RZ�v�h^�Y��7���Ƨ>�s��;6� ��+�wY�ތ��t߷ծEU��Ã~�+�L���rK�ow�L�.ps��#}�)_� d�{{4�O7*ᑧ�@�5��S�'��(���or���M�q�3.B]�wm��s8�}�s!1t�s^Q 3�$ֽE�[��ؼG�[�嫕��L��36;O<��iy��'/�����9�q|�]8u*2���u�}�i+}��e�]��O��DC|��Y��.웱��V���k!��;�e��i�$g������/�\f,+��G(���%����3z����"�"38�VN�l�P�&N��F	�`4�M��:^Q�#/"�k c�Hf������w�Y��r����Z����ONeq�ۇoo\{�}�.�M�^�#5n�CŹc������p[����և�NSQ;|1'�ӻz.����{w��!�֬M����f�#�c�E�ӏ"�{������qN��������dW�#G*7x$;a�o]�å�g2�N,b�1�S��ؚ�X�.�<�u�>wQ��g��s��^(�?���/�N�S.�׮vy����wY����k;�3L�NLw������Zܭ��熆�����p)��&h��M���[�f�4��?g��=��{�>G��M�m�/>�g�����3�b^C=;*��Ւ�堏u��qz����K�B^xv':���]cR���@t�/���7b��S��ş��(��_k�E⏬�׵Ӛ�{��|;4�f[�w��tנ˕��M����_�p���b��w�#F�9yD<�/��;z[����2 )�m�;��onum�ö�UA����w� ����=��X3�������������9"g���΍������2�x�=�}�Q���ۛj�z]@���c��a����'��dβ����9��bOPO��a�w�Iv�=����zq���S�`�rM�}�r���ު���u��:y��w,� 3�}��k4���l,�gx�K��8x��� �{���w�v�;�D˪zgd�9�ӮA&]P��wc��^^�#w�Uy]���[u����A��r��r�^�{��[6�x��WG���� ����l����� s�/�b�œ�[����m���Pz��9���:����&k�hu����!��?:7���LY��,�9���FQ��o+F�R9��["�����1�q���Cy>>]L`�x�ޭ�Zq��/�h�H���%�*�^x�W§ΌWKͺ���}�gV��i�y�9MU�:�k���NTLO��{��t���,C�n��'{���Sv��kN��t�rn���ٌ����9v����^�[��eԜ��":�(�8m�njƪWyL;�c�}�<C�{l�z;�+��ӏcv��/y���8Ь[J�o����U!�n%�v�MeT��yP.w0@z��36e��I($M��1:���R=�n�m����Ƶ,���!{���2�/��!����=�*/��9�::��Q�K��ӡxY�l�[����{���`:w��N���)����wڸ�}�Y���JM���\�"�io�����4�T����<�I7�̡�{Dѓj7�hqr��D��du�46��_w�<�g(ʢ�E$l���;&��&�ɩ^R�sL`N�w��it��K�s���;E-۝U6�C%`ңq�Li��AF���j�I��n��53^��,<۹j#}6;P}���Ɵ`�ٳ#y���V��ցۆHܡ7;/<�8��=�Fn:w�1���.4��T��-L��KH��C(�:�*00�̧Fɩ�8�f8
,�f�9b7�����OQ���vT__?Lz������|{��[V����N�{��7.��ڡ���-�1�vI��蓅k��
����G ̙�f��ώ�께���p�Q�g���0���]l`�.kfvu�Z+�F�A�z���9�g����
��/4�c�CON���I5���b�wܒ I�G�%�|ܮ��]X�xW��{�+��
K��)��.ZX��sð 5�)9.Ü�m���A|�~���?u�J�e����;p��7O��0.�lX�l!s��=��{��\��5[�t�N~��M>���٤�)��ަ��9�_g?{h�{��3��Z/���\��]��x�!K�}���$��O@n����}3�;�WC�#ƃn=�9�T<+�''��p���졕Q]='��d���<�o��o�l��ƙy��,�}� ŵ�q����� �.��}v�}��,����v�w���nv�ո{�>E�Ve�f����/,*���n��b2Պ.X������Dz"$������?����O�~?O���O��h�5Y�Q����-�\�S�^����a���S��%�㶭wJv4��1��i8�97�YL��Al�nu�fu�.6���zB5������4��n�t=��n룎.܅ tr�Xs��<��rv9�룷k�t�W�SMۛn1���9�W����u��.��'h�^�^9�ض�w.�p�m��乛���ې����\MW/U.c�[�(�۴�\Du�[a�靶�Gkg��i�ӳ�b�^n�%��u9�Ë.�[u��S��3ױ��W�<��晎�k�؍MS��z��4y&j��*������|�;Y޺7W3����aŭ�=����=���ާV��������;-�uɬnw�z� ���B�yc�$�v�`��/���r�cdy�^����\�N�N�m����ll�.̅�sgY�b�1�ۜc�v�E�=N�Da�Y��S���E	+��p+�u�&�p�q���W9��r�4\8㗶U�����ť��]nH���`��ص�۫��vk��7T�C��+��pݽ�ڨ'G>N��s�\�����j6�u�9�b�l\�7]��۞z�o>�-��kn��7QE�F�!��I���c3�g��p���uՎ6��S=��n,¾gwm�m���Wװ��"��=�ۮ^����U�lv��i<� ]����&���`���do'�k�d/'�zI��9�N�n��*L�,K��Fu]��]�Kx����!�g�\^�郮�{v��<t#���u�n��x��;�n��ݝ���竚&N��r�H��vP�ħh�x�]���V3ť9�V�l�g�0��=�nǋu�өt��Z�9��\�i��Qt�v9��>=�mb�Ã�X���vq�-��Wl=��`��n|Fw�3���y6r;��B�^9SŶ���.9��@q>���cu��^�Ѹ���c�X����e�Gh�o
���)�P."`�������kqZ�Wm��;<v1�Rڛ�n�nn{Z)��GZ���c��D(`)��3��Q_꟩g��t�٘�31Z�$v�<F+iz�Mj��T����{7@��c���_n��}�D6�Fh6%�jo`����6�+@wٴ�)�� ľ�U�Y�n�Sޓ���z7�W��e��'}����rg���J<��"��
n���������}��懋�����>;G{�ʹ��g{S4���.&��*�����Lɩ����1(3K�v�6��' ��:�o`˗!�|.�vmZ3��P��8��J=�0~[z��;v
�/	t�53�&è{�F}��k���Ѻ�Y�-3bspS��ؽW�+	&�A��7yo䡆����Ns���77�pI���y��=�Z1��y�T
kf�Cz+ �}`;�'[%�B[�cI����x�M�N'�7�_,}��y�5��������6�㜶d�&�s(@�G�'�����-�h�d�鎓������[8C�og�J�1��*3�*�����=&l�(���rF��l�UVE~��KN[��`�M�4#C�-bQ��bUd�BV�ḭ>�&�N�pæ5�9[O��u̻������V��<d8pxW�D� d*$�O���zֽ�ĺi�����UY����l"�O��o/
-#;�T�\���k��{0F�3��<7���s-w=�
��S"�@�v�g���c8v���>-]�,2�����Y�G.h.ji��2nvA���ԏ/,�E���V��%�8	�	":�6\�F͉F�u����8nͳ��| l�E��jwn�od�\���u��G�k]� ��uͧ���B#v�=���㴒���)��]/]��<�'���o2�ǹ��Wn�����λZ��s�	��:q f)�:��u����^��;r��=��y륣�^�pf��>��a�.v�9Is�÷�$��Y:��·�=�g��Q�t���.�\��br�g:9�w����ѷ.[��.�`�ݠ�4A$�Ys-�M�2Ph2�<9Ȼs�����w�cm�vy�l(�v��R�N����}��@����f}eoWጶ�Q̭�An�8��RF5��������f��I�M�إN ��ð���8���jh�T��a�%��3��̑��f.���S�����`��~H,J�މ����&��[wJ��u��/�\+�o��	������v�͕R����߮ݼ.@���c��{�" F�&��� Ц�-���x�`�wN�z	��O'8z��f7g\�՗�d�3X/~������(��q-\3ٙ�H�^f3��,��a�CE�$�]�x\�'�ǣ㉊ر&��<���fnw��Z����v�kt�6���5,��U�g����x(ݷ4��=8{��h��̊׷�����	�+��qι\�;�r�)wk�Nw;���]��r�3$c�s�;���Z����S4I��Z��!ahXPIB�KW�2��k1��>�9�߮�=.@���q�e����"Q��fg���Sb���E=�a�{�/�!m-��hX�B�N�c1_�H��}���`�%��o�v���2.Я��w7$4Ԉ���LɌ�G��]���K�iW��s�\�M��=u��k��]�ZD��1c�T*�l�*e�w+��[�o�5��2��d2�B ��M��:����+2yTp�T��L�7baOd�p3�0�%	#wZ}�LʭG"��u<��e\��C������؂f��g�=m�0�J�k(���\�-|9���]��͌���r�na;�E��F�,«�βrtFauk�=��긘�ۺO��t��x��-;����[�r9t��(E���9���ȹz�{{�΃�.�0$�D���}�?�d���&"Z��[�ϙ}���C;ι@�P8�l"R�f�Ā�o�*�,��5Lp�4��L�}���~~�.���۬z��s�0Y��x1k�M�(k�4��Qf��UZ
�v�Qu-\1�֫Y��|v}���_���i?Se�1#R4pǻ��8�������*Z�
��.�Nz<����@iH$7�(���v}"��c�+cީ�=�VM!�1¦������'���� ��={����sv�,ꥸ{�`UF�X��'�!;�^v�
w�,�NB��e�1P�H��b��v�r�҃/(h�3�B.vjD�Q�3�'^}˾m��b�* ��Y���]ݹ��]�wr��`,&s��wq�9a�f�_>��jW^Q����P��"a�T��Ҫiw���Q���r��)e�U'}�O=�m�N�;E�\"�9��l�oj��c<+o0��������pU��o������%��V�Dz*�=�S����P�&�M�� ����}��Ktj�6VQ_>�g �@Mo���
х�j �^�kzd@� �O}���(ʽSeV�'��Y12$�y� C��Y��i^#>�;�D=�DR��$�p�m�1��Pǜ͜�ʵoV�`ŏ{Â�ټ�Ne,/�F�W�3�[=�mq��W���Gl�n�ʌY�&qWW @[�fe�p�]@k�9�<���'���]D�Z̜����Qia5zK2YC���z�h뭂�Y�mԘ����f�ٵ��l۪�[N���K��xƸ��g�'/e��ح�֮^�w0����G;���=Xƃ
㷴� j�㋧E`��y;l7��"��lj�N׎!Mۙ�mv���:#wR�<�aMq�g��+��z�]i踫�Ǥ�w=kX�ù;q��\Y��>qg9����"NP��վ�+��d&�����AQR#�oËŹW5���(��5͹��$����Rnm�~w���~Q���j��b2���v��X==q��H�n��s<+��z�D&�ifQ��>�*����_Dz�2t���,=@-�m��!��V��	�~��-o���d[潱���I��r
�5����`4@3m���Y���1�u�qwH���2k#3	�	� �i�)W{�:���[�O�J���;舙S�5dݷ��L�	@`&D���b�ߕ�MW>�{�ᶥ��d2-���>_rgTP"LZh9H ���f���[θ�7�=n.�=�1���/8�%CL�w��Xa��!���6"���*���]r�c�{ǃ1��þ�#E$$'m����������d��ԷW�5Qf.M^3�=y�o(�E.A�gPSoE<r1F*���aqꙨ䷤]޷e����^�:��5]WUC�d�w\�w\wq;�X��y�H��4�HEi\Ws�.d�X�H���n�gي7���I��B+sQ!�^��zZ�fH}�}Z��M��z"T�x���`����(��<�X�R�y0ęH�u5��z��JRѬ_$��6��{xp<̓�	 ���m[�E�H�H�����A���QB��v�.y���V:M���0��\]F�s��s	l��5�0Zz������T�p�sv���.�Tt{�v�Wh�UT���5��I�
-��v.\7ڠ.G�E�E7�=d�r����W�ԓ��p�h�_��yʢ�S0T*�@�gOr��{V%�I!E���}��٭�7��ȸT�	z�%��b�uY�41��ki��d�q#��s�1�v*i�c���9�������|,DwtbBD��w�]ws���������K���v)����bZ�q�`���^I�,4A�n�"=;UM)m�Ѯ��b�I��y�)���~��4��Ӆ�$,1ĩ|2����H������g�/���
.$��m0�*��5����U�j������@.+�M���v����}�K��l�p�}����xf��n��D8bD4��5�D�gb=/�"e$�F�U������\��0�m�� �"���Tl�z""Uf�FVc7V�9�6�D�h�
0��
�"��ii�S�{,I��[̌�[W"��\+�۩N��p&�n�H��d!1Ց����D���ʪ#.���u�q��r�s�B�q���f_FR[K�����T0်L9�bAHa�����i�˻�s%�[\���?��40�� ����C��&Wz"3�R�oe#�����G�_��G����A`B��n6�nϨi�݊��a��*����0�us8�fn��u�%Υ�T��A� �c���Ͼ�+�ݷ��HaDa�0d���Z��pPU��S��}/j����
���hԱ(�c��xc,��^�32.�%c��?��e�#C-��1���&MlDy��[�ܦ$�
�b�����:"�����eCaC$(a�M�4��J�����xiRF�M,=��t�e
R"՞ܢ�U�6�tReP.�О���;�wu�܊��|o��޼��0,�ItB�|�G���;7)�s~���.X����ϱ���0��0���8�8W��7V��:�jv�7���{�z�q¢�7Y�y]���8�yۃv�!.��
��Bl[]�\����kAf�<�gT��ݹyO�v�9 V��	�]���w9��q���v�N��g��ֻ�A��v�����m8&�cp�\��g����I�F�,қ2K�>���t�u���܎��Z�����h�Ҹk� 	�T�F�%R\�+��:
r껻��I�R(EBW,�K*� ��A�\������}g;�Y��z�m�M&ǷW�ib�A~	��m�I8�-�r��e��R��?{ԩ�!>�+wh�0C� (Af�$o9�Dz*ޞ��:]�bL����� l�{�"D��4T��Ǉ��Y���>ϲ*��'oyG~>�� h�`�ƊnVL誝����p��ҳ��c�w;&����$��	8%��!z�+h`�+}�5y��֞��:[�E�}h���c��!C��q8�nFTREA�3ds�#�6�$��݆%)7U�"�Y%Ba��d����S�dʻF��&�~6��:�,F��Sa��T���^����U'LM����"6HQs<��"�T�U�z�{"���uWSy��hB�%6����@TtgA�N�����S��j'Q;@�=�I����2ή!��٨�Ĉ&��AQ���=��|�������1cu"�l�P�$��[�O�J���[��Ӛ��-=��t��(Z!�-��6�tz!��9\����S�d�PΌkk]���>܎E h�,ҥ��SK��]��v��uE*Af�U8�B����������q�#q9��
;mdˮ��Ȯ�x�F��]�浘[�S��	�k���V��un�Ft��72^-U4�G�Y&E�N��-���y�xr����%J����Щ�yɒ8�X2_�Rƴʕ���S~��7������1Vc��8�2ތ�P��e4Fu]���{���v�#;o�����c��x�}�o�q�P鉙̶0��"LÃ���+)�svwS��9��r���z�zC�h橇vln�e2�=B�E�V	f���v��O^Sٱ���'�N&�jo�Ĥ�3L��ދ5�cUnDw�'!��']:N���:P\� ��Ыq4�n��;˸"��$Ywoh�3͎�qi�]�Σˎ�$�[�/�0{H�NR���sڶ��S�qTH��7i���T��:4)ݯS��h8iLꃺ�2-�n������N:[�i;XL8�u�2��m�|	����)��v�������:�r��4>)��� �MM�2���(�}6��A����=A��;�9�㿫�k��ܡ7��|�b�XtW��sn�n^fFQ����VS�鑡o4:�
P��t������K�;�w�z�Ğ^MW���g/M���7��Z�>��\/�F�~e?qC}Y���i�8�l��,^ef�2T�bF:���M澾y��1kSR��Y���_R��R�cMWq�1B�q�s|��S6#��ʥ�l���b�����;�����Ol�ub���_{�X}�=����s��w�reE_�x)�\؀��,�7�ܣ{���߬�4��-��� ji�L�Y��S��j�@1��c�kֶ����XT�b�`5gu x8��Y��¨KG㻑}�>=�u�gvЌ\P'S�;m<��,�K�N{@ߨ<���F�}��0 �;���t�����������q5�1t/g(��crU����(�uT����������o�A�{�Λ_'�ޓ���7Q�1��Z��BZ5v��x�[�n,cv�I��l�ZY ���0Ue�~t�d6V��S�Y��cNa�*��I0DQ[�qJ��li�bȽ��D)�a 1� JFљ�]Z��D�:�X,J�\�,Z�RL�LAY��N\f��e��mr����Di5N��Pna����r��1���k($�J�B��Ұ��lҊ��g��;Z��E�%/�g��pg�9�p4�V����Sg������U�͜UG$^���:3��p��#�n^ѵ�*/Tg�-����P�70NF�l`�v�.�ς^�����i��Y�B���c�; /��KY=����{����X��6��e��{�V�4Pԁ2F-^bʇ5k6�ɳZ�s��`I%U�eυ�ұ�47E �kҜN���ͱca���c}!�]٠e��WnLڙכ��4'x��p����S���H��EanٌؐmA@, �k՞�%�tW\K��r���� ��z �Ę��sc	d��s@Os�Al4ેC�L��/�`m�8���\p2�K�X�&X�����$�����Zu�y�1� �wv�''�w~��燞�<�`��7.��식�:�X�ۻ��vq�>{\��G8F(.�1���6�g���Y�Zm����카�m)���v�U��j���$Q��XF�@������#4��_oi�M2�|�jT�S4�f���MB0�!O���dl�c�#��H�ZD5���X�/g�T�^�p�y���{:��e'��i)�Jg���L~׿K��7#p�>��Kr\A��g���L�1O[��.�Ԇ=�0;��P�-*A$_c#�P�v,�XD9mϔjb��o��6x# �m�Kǻ���{e%}Ю��rjFn�"�"��u���A��q��ϷSIL�S9}�Q�gU�5�|��U����Y��`i�<~S��/��8r�P }~�~�|�N�<�~�;h� Qp*B���h��
 _3ص[���o ح\ǰ��u@��o>�r�ۢ�n�ebا@�0��+v��%�i�4Bx�1	�1�;!dNi���Ud���,��yW�������W/����^߄�D)�rH�����6/
y�.qݮ�\D���>gW�o�ٍ�EE��[��|�>`Ǐ��+� �侟>�]�oZ�>
�?���Y�HS�B[j"��ɩ�8��ڸ�n���z����5p���V�G�����2SPBp�L�^ŋ\|̙C�U4Ͼ����@��~�~��犃��E0�r&�yx�\���
���;�#*8����C�T��.�%$T�b��76E����ݝ�}ѻ<(W�}�~U�o��T�cI�6Z�Y�l��P ����O�p�fC�����誺��o������8��aע�H[e�ݛ�^�!������5�CZe3���fY�Rs�jT�2�%37������ÎN�(
���^�\����V�#O�Դ�*��)k��K��,Z�Bm�:����'��K!۹���ȝr�F?��yY���H5��5,C�q	qc]/`}���rF�w.��`�N��`��9]�׳kV��.��{oc��;n˞ &7<��͵r��nwT{X�������G\��"yb�6��$n��b�.2p7�3�;Q���T����{q��R�vz�6�=/�}�}�s�ۅ����s�Lt�-��[vql�nK6Wn�n}l��׺vݛ������O���w\���sw9(�;��5��U�QIwF"��hFd��NCl���E�-,�ǣ=	����^9�!k���y�qɶ+������۾*.7a B7_�>5\�/ˆ��5�����:ٶi�e'~�u��"ȀN2���4��|�����>yQ�0HVk%^��m��_oi�A���I�ƭ(�e�Y�fi�M0{\��I���
��kg����FbQ� �ͳL�)9�^��q��%3��ͳI�N2ӹ���6��2����3-a�B���H�K��A$��՚ސ0 ϵ���6��m�u�;t�&��S;�{r�x6�$a ��o~nq�ͤ5��F�$eC#�!��Maj����4��/������6�l�}�t�Y�!�ݟ)Xj�� ��8�%9����m!۴��r�lk�m�ڵ�K�����L�[�ݯ��w�����թI*�j�tͦ�e���ܳi6̧~��șm)��|�6p�I�m8�N��V����58OWpDą��2�EcM3Zj��X[�{����0y��4�$}�t���`or�w���y{���w�D�1{"%�� 7wmڧ��J.��m9]Y�p�W�]�j�K���c�Uc=1��$�X)g���r�v�Y���%3��`��Ri������6�f�L�=ΑcMx ��5�7΋~AG�(��;�iҞ���Xt�G��kU�!�[9��(�2�2��L�3F��k�� �P���2�Zj��-3~��q4Ͳ���^K6�I���k�ͤ�x	!Lϼ{w>f�f���Qp*B�ѭ"�P�_oi�f�O��0�@'zrfq�g���pT�)4�Jϸ�vͦ��S:N�~?7�^{�,Z�x�稝�Nc����O]�Se.sQ���V#���u��^z��1F�I7*�Ƭ�ơ���5i�;ӻ�i��)>���<d��[6����,�P�wJ�dQF��
��ճiL���SOH
 ��e��=�f�Iǌ�w>�%�e�l��k^nm=@P�_f��*Ǆ	��a��(Isl�m������Jf�L��x�L����>��a}���}�T* ���2�>b�+��t�$�UcI��I�S���#V�̝蛞F^��R�㠫3vmu�-K^(��G6'z�OFdoh��@#srr�!��ם�P��A"BHQ�
N�\5���k�ȳL��us�)"��
&e�il�a�@�}��6�I���כ�I��1ޝՒ�I�F);^�ҙ���;�\dC#�RQX�L� B9�r��RJz`��捡I�RV}�ڰ�i�JC����m��B��6�����m�	�1�=8T�䍙��j�c	��ql����m��)��f�׻���h|��p��1�u�!�CK��Ei�Gl�e��C_}tx�$�ٔ�O��r��L�����#2a afƑZi����p�����e����i6̧}W�ɖi2ϳޝ���A$���+�|@`�$rK&��kơ�{,���4�Nr�J�e'@�@�[9�~jm��e%g��.ٴ�6�ex��(d�#Q9V4՚��B��|nq�ͥ2����f�l��=�,�S��}e�C��>,����C���h��ޒ��!�"nM-����TeP���PA�F�]����]���u�V.��ݎ;4w�qW�v�,!xI��$�"&9�A͊4X����@�.r���mzo>/�"��!?��T%B�JTFF��,�e��?54�M2�� ��.���8�gs�nY�[6�O�Z�si��ĳP ;3��"CI��Ka�*"����K���d7T;A#p��0�$$q��� ܵj2%eC#���K��ϔ#��	�%&��ڷZ�4�Nr�J;��l�,���5�P��x�㑒��`�g5��m4Ͳ��k�䳎�	�q���o�Ͳ���V~��UͳI�R}��&��UQ*�֚�W��;�&$Iā����l�2Ͳ���R��L�S7��SL��m���w��gL�)�Ͻ�cMY�5���q�R8�nCu�S7�b@�˯��s��m������%3L�o�[F��i: �!i���fٳY{�XA0�!)(iCu��j���.���6�|`C��rr�q���k�ͥ!��Vyޘ��q�N2�ﾾ/؈��ٴ������'���Q2�@����x�nJ8up�Y��y,�!f>�'tX뺈'�u�"X��`��̋�U��r{f�_C������>P���8�������ͪ�6�'i��H��j��������ܨ�8���m�k�#m�6�s��e���z���x��)c^#:ͼ.z�[q��'�<�Ǆ �wd쐯V����Y�q���}�~�lv�=��A^ӾnZθΓ��I��a���q�s��B&�D�.a�Ò��#�=��f|$P���-��X�L�-����)ur����<{��m˅D�s�{.cCöݎ����ww���x�F��Ǡz��cl��D��ɸ[��~������l��h��D�!?��(�6.F	N�(	rѯ���)�~��3,�)9�S3L�4�������0��-6�LW{�]<N&��[;�z��đ7"3Mʱ��֚�w�<���FHKg�y��qW6�&�I�߫�S4�f�մi��!	L�->=ߊ�Y��Á��Uu��֑q�L�5I�Rb���]3i��" Kgs�rY�Zm���k�ͥ!��W{�Yҩ�Yq�4�UT��M��	��y��S4��;�h�2�B��534�CI��UB�}3� B0�#�<��$TqSA�ԉ�F�!��ڱ��� C�A��~nq)%2��|��M5㾘a��>:���0��<��UņٝЋ�ծ�ωv����d��hmi��  +0]��H�mT6>4����534�CIL��ɦi4�LW���Č���q-�Ͻ�f�i�Rb��y,0Ϛ�£HG֑i�s�K*�������57�13����j�\�;=��n'�NA,;ȼ�7�#S�)\eut���3]����Q]i.�X�=l��ǭ똵M���f<"�� x09��.sE���ܲ^.`"*��0�zI �a�&��54��2����4̳L��L�'�D� �ZE�Vyҩ�3Q�R�5�i���{غf�L�)�g�ܳi~��C�Y��u�kH�Nw�;��=~���D��R�$q�F�0��
P� Y�{q�l�4�O�534�3IL�o�M2�I�A ��7��L�sx�e��W��qCY�s��f�l�);����L�S�3{���3I�Rw7��4��5o2���v�}=��� ʀ��/]p�;�6�ے�-��{$S.:p��V��z�i'�8Ur[T)D�JTFF%]|t���t��0�!N���#i�x�ݫ 28�3���כ6�fҒ����2�q��n'u�aj�}��d[6�g;�h�2�%}񩫚f�w�#M*�Udi�!X�./F�rC@cq\5�a�5u��V4���bxS��C:5��F|��s@��\�هћ�Y|b�p�b{bgnQ}s�Q�������ځ����P���B�L�i�N7�����ӗ���Q� B|	#3D!`��[��#"W� F�b>T#>���noK嫍����Zp�]6�w|*�
;ѕ2���fL|�ə� AUBw�����|��(�Dc�����y�u-��PU��Y�ά�g���|�>=�R$�J���,ty0Q�<�4��iy�Yt��u�c�"��Y�߻���b
(�)O����f7�w�[ﾝ�y�� a�{�s}�fD	N�(	bb���ug����82�[ߚ�f�q��U!T�s�l0�eȁlēpn�x���Z��
�*�}�a�IS�4��S�d����F���U1@�mh��gz�nl�9�ڱ���s��!�<{լ!��Y���:��7u9���)t�@0�0ܟ�;��~�&7rnB�.�/+���fL�]���=�=�� ����z�����4�����]v%��u�		3��}�m������5i��V4H�r�����޷Tc�2�ҙl�Љf��(�-�e&9�R��l�S7�Ff���m��g��?�����sX#�k�+�$<W^��v��ں�삚��O
K?��w��7�V��q���f�M3��w���6̳l���k�Ͳ���c��`��@8ͧi��dՑY�k�x9��ȆF#h���l�m���J�{$I �6��|���4�e&=}�n���6�g�z�,�= UU|j�V|�J3�q(��u��m)��t�M2�L��,ʗ]�f2ً�أl�i��xԳL�i)��}pe�����Wp��f�od�-3�{ٺgL�)��rͳ,�)>�k�Ͳ���F@��=�ԩ�Zi����9q8p$hY5�CZj�樓e3L�D����M����sՍ4�M2�����6�f�L̜��ouz9������=eP�]��a��c�{+�2���x�n޳C��8�=�N��aBq�&��pMV��ѭV�\�r6�C+�:O���n?A��]>�����nپ�{זN$�C��x��7��a��qT_�dJF`Ҫ�d��z�Q�: �r������1#�`nzv�>������G�=1���%��gz�`�ǣ}҄H�>���Q�M�=3)����Uˉ:���Ŋ��� 
@�~R����wzmk�1�������oWOkB�-��s�B��ُ$S��b��}:)��]V��U�]�E��`�빡P`#6w�K�g:E�z�8�����s[�R��Ď{�Վ��@����s���dc�K��!���o�����|�䫼�;'��t��_~�_�^��9�M��'�P3����N��F�[�b�E��Oz<���E;.��I*������Z�"2�j�J�5L����R�p��X=q�5��� `�wo����݈I���l��/���.���[�m�Y��6�B�}DXs"��1e�[I��-���9&�u��V��[��ΗPwvc*��w���y�\[�ڻ����8���B*��kp<�Ncv�k��F4a�Ij@`�s\�/�v[������܈M��?t�6�~��ãx{�3���4fފ�r��ޫ��VmfH�f&/.��:�@�1���u��"�U�lP�"����2Dx����]+7����8U&�A���=���޽�|+K~	�8����7��9b{GgG`�{��>UGM��/H�������y̽��iv�W��٧d�v�~^�Nq�u_E锣�<8;�$�@�2Q �
AE6�bf�l���6����EMn^p���Ȁ�1�c�R�&��7�_q����ƚ̠8�[��ܨۙ�7��u�v;kl����u�g�\L��	$�v�B��]U�e�8X��[��n�������^ �bI�3F/n�-g���&���ì�J���59Jb*5��<;�����,p��/]g��g�
�nq�cq�W ,f�r{yn,��y�X�vμ��_]]�ɠ��3yQ5qՎ6�0��h딳;e-�p�w"������z�f�vչ�<m8�4s�4d6��Wm��8��>n0S�W<�cN땸�'�v�A�(���;b{l�g�ٌ=����<�D��ԛ��0e�N��r�Sh��^7<mmWlu��q��wl�����.�7`�ٯ=����ɶ��gM.��lr\�˺����Q���֍�ͻj�Wqy�;�)^�76��0s�γdv¥�m��u�VՎK���p���c�=�;uEç��ţn��N# ��3�ϧ�v�[<�n�a�z�y��3�zC�w==���n����v<m�2	���&;;�;���{/[۬�z��/
�fY\]tvj�y:�1�,Ӊ{qva�E�n��OUi={F��ι����oC����O>��qF��^0�/d��7n9�����[g^wJ�G�@�'��r�l�^��j��ɮ��D�'���-�ӎhU���]�u>-�{v��s�po[�ǐ2��T\�ѵ�����꣗yx.��x��C=���p1�e�+m�.�ú�^���]��Ƿn�����n̦�]:j66����.,�m���=b��1��!��bV���k�0��3�!g��ݽ�s�;l�A]#W	\:�ۛg�*'=�[��'p.9�wB���k���Ogr�m�Oz)�d�/Y۬��[�>��k���n�x���&['�\]�,�J\[��u۵���ݹl(4y:�/n���T#s�x����2*�d-o]r�N]v�ͣ��*��<��\m���ӸM����p��n�I3�:��}�d(Qq�78^z�	s=vN�݆2�K1�g�sL�3�L�~�ʩӝ��"���_��ˬ�7&���"f��넺�7����5�7�:=�G*x#<�Jqf����_LHvQv���N��r�T���%ѿr8���u/]�������i�-ҏ�o{�����T>t�d��c�Fo�CY�b�&JS��q9��x}�pQ�-7 GǷ���Nr�_+���W^ʃ�����E䳰�A2���n�8�TP�0oU<��-@���m�5���hDC���[�9����⛞�y�t��as3�xSm�Z��"���af�FC����M��2���A��i����1�Ԧ3�j��=��p5جy�R��������� �$y�tf�F���E��5~q�\�AС�+0ƜmS�4��x���pz���g8������uO��^�E�d5�̃Ҭ��}��~#welkҨ��X��t�2�p��g�{�h!��`�zfĊ���g��<��-�������ܞK=��gB����m{����Qp�y�+�y? ��+f� ��<�ɸW�ok{���(��_���'�P�>߀޽��w�l~��N4)կo���T�Y,u���+���n��Sh��X��}�V�T��rN�r�Q�|����{���� 7����W�������܍����I0oD������4w��;�u��΂��$��һ�&���u��v�k�&u-����=s�0Y��ݛns��΅�n���,b��ݝ�q��N��Ͼ�|�T��a+�ms����1�f��;'�_}�l�n ,7q�F�']�4�!M�ǧ�f{0���f�Q�u�W]��7m���ݹ�B=Sz9bɱ�k{v��.+۶է���۳9��r
�Wk�$2��>;��wPnWh���kDhБRTQ;��z�Z��K���O#x�s����V+ڧ�M�vv�u���Z�V޸[)��w��{��`�L��-IV0�5�P�zg�֚���is�R��i�Rc�h�? �i�m�Ҝ,Y�j�B��j�)*#!bK�e3iO=X�Z��-6�Lw]�n���6�N���oFY�R}��[�OC�QV�k��G�Ȕa��Hs	sl�m���R�%�L�b�r[)� � �-9��6�f����*i�F�(5��Q��'Q�p֑���!-�ﹴ���6�N�����L�S1����٤�x �	i��e,�,�����}���.�CcMY�����jT�)�JzH��}��6�M����7L�i�e3ｽ%�fY�Rx
�x�N8� ���c��L0�sp��"��h�Z8���^y����I��/.YF#��|j��iw��E֚�4�!v�YiL�S1��i1C�6��T����k��,1�jQ��P]i�F��.ߺ���n��ľ<��K�k��ڞ�T�������F�__%<����7��|�,˹v4�ͦA�P�		��%�;�*��챗ݼwkL����\�>���}����Qb��CƮ!$��e���������nr�\g�H,�e���Ifٖm�������L�S1���������m8�Ow��2 Jp��R�Mi֚��l1l�[)7���4�O�����%i�F�.�z��0֚����l6�%ȉlĔ��i����� �k�nq�ͥ3ﷄ��i6�Lv̬��Zx
d�	�\�&�L�Rx���r TP'h:��P֑{�`���4�{$@!���l8�g��}�%�fShRs���6��ҙ�6���q��*m��wM�cY �ݴ�c�볒6N(��v���-�7�y�߮��q�@��[�.�a,�'̤Ǯd-)���7fKe%�I��ԣ�KCil�Սi���K�"E�#A�`if�L��oIf�I$)�e�{[�sl�m)�ｵ.m�M���+-<H��,��\���FD1CE$li�kMB<�2�a�k���X%a�9U�����ٚ�n/1�e��l73�8��J*�gr�(F��zo�;�CP�LIػ�]T�. ��eWd.]Q�/eGv�Dt�ڧ;���7�sWʩ�A�Ab�V"���#��0�C2&���r.�����Lw]wtͦ��S=�nQ�m�e&)�r,>� d�[�Z|E���f�*��W}�)s��m����YiL�S1[r[)���� @-=|36̲�=k�zdhD�H����$5�=$��wR�3l�)=���m�ͥ3w�H��#MB=B�=�,����1M�k�:�zK�ނr��Gbu��qp��u@���7&V (
�nN:P$�H&�X&P�{�T)-�3��M%!��qe�!	&���-1]��l�q6�%���<��E�V4��G�=��} 0���[1�{�Y�4�e&=s!iL��1[�(�> �@��hB��=D�eFdhʺ�!H����iM2�_q�U�gi�>I�@!�4��(�6��׷sl�m)�_os���F*�`�+J\�4���H'=�+4��^y�*�fSۧ�4�f����X�����vi��N�g�߭7w����n���Z&�$�w�O�ftH��QL>���Mp(�˻=;��,�,m�tIs��x��� �,c��&�Bk{uvf1P%lJ��Jd�e&H@���54�a����v5l�Bp�ikMC_r{j��L�)��$ݽ���S8��w�ڗ6�&�I�ٕ���e3����w�ߪ�ٝԘZS����zv{��&�6��8Kb�ݧ�7�ww{���}���r��UX���q���:�4�f���똩�Ri���q��= �I'l�-�v{jƚ�i;�O��#A�ገ�76��ғ�{�qK8��H`		���L{s!iL��1���L��)>�:�4�Ba1 H[6���ƚ��W53FC�����j����0֑>����C�"!�Z{տ78�s���S[��Rs�W�DHNQJT�ɭ"�
�@
�!�<v^N��Fh�򕆡G �UUB�w��\5�kMC\����e�"�IIV4�5���Λ�5i�����8�'I�Y��YL�1�`qC�=C�AR+w�N	������L��r�U%=r�鸾گ&�v�vk&�3��d��6��%bP�y�	�aeJ�5� r� �{�:v��Ka4�+�>��f�l]��5d�'{m�W\��v��.N�z�K9���FvHJ�;��8�W�ܝXT��s��q��Y�g�7n��C���]��v�Oa^��U�r[��W�֬t�mf�n{O��Sm��.g;�-MѠ��㷲T{s�T��'A������J��p�������r]���<d�5��ŎD.]�y�NS^�x��ь�ɸ.��}5>�60&�߸�4^*�y�E��Rf%��mK"c%�`�R#!�u�`�Vk5�%)Uի���^)+��{zgn�����[�烮�2M8�A�(P'vY�Lj��WXj�!��e�Xi���
s�N�H�ZD5�N�Y�H�i�Zwժ�L�IL��hsԄ�7E��"ƚ�4�!r遽�����l�)���F�l����Ke4���� *�(l��S�2PN �b�Y/�g�5��C�Vi�� ��)�_ə�|�e&>�+-)��f��s�e8��6�P��P֞P �����Sl�i)��oi�M2����6�|�BI�z�ܖq�Ͳ�{�1�����P��5i�/�:�XF�ċ �FVi)�e:L��e3B9�9R��5�C_ �<�m����^36�6�3��v���6��l���R�5A��u�( C�Xf̍�H��W_i�Rb���L�i�e3�Ww,�)�e';N���Cl�m-��XL�3I�R89�%d4�I��M!d֘F���@[�m}�іX�����]<7���H9����zW�?1,�����Ou�>�S���}qK�K-��dZY�0����GH+V��W�[��ٷcrx�� � ���d�kQ����6�`�*,3h�4X�ɢ�F�X0#(���ĒfY��XJ�e3IO���T�2�e&+�{tͧ`�@�@i��Y��P�C H�14\rY��o/���ٹ�[6�ϻ�&f����i�{��m)�e3`�e��!L!ti�H�PH�D]i�k~ �I�HC�]5Sl�i����l4�a�=ϻ�f�I�x�d�!$����=��"�D5����Ȁ�M@L�DE�!i�R}��L��=� 3e��g�"3&O��,�L�5��.u���mp^�׳�6g���N�5덮�]�{R��q�k����W�������w۾�����J�M'�kۛ�L�)9�^;��e�iO>�'��I �6�KO�fVZe��4�x�|���al�౤3���a(:`��%<��ֱ��Ϻ��M$�=ϻ�f��I	8�J���f0�-��CZD5��!��0y��0��B�dN�d��fQ�3���}�&�a�G�J6{��
H1��o*]��Wf��{(��X4v�>ɉ��Gـ��ņ�ݠ�:���IZd�/�W"*$�9����		$�,b��Dst�Q���J#Es�F�)"(��I��,�)�e2��������"���d�Lf(������ٔ��A�����Ϯ���m��v��f�L�)9�_qsl�m< ��f��D1���5��W�DHNQJs,6�fҐ�)�JB��2 k���ZD i�/��@da�B���4�5�Bht�]���@�i��7"c��v4�ۧn�M�K��N�HӇ���W������A�#iD��%%X��#�#���.m)�3�k	�Hi4�Ng�J����m-�l�]��=��3Y��NisXg	siHm)���4� 0���-1}�q�����=���e&Ф���������Ķ{�l}X���R�a$E֚�4�#��!5�CXj��f^�$L��+xJ�e3IL��^*��#B'�*��%�R+���3}�b [=�rQ�q�e'}��,�[��"*���X�~�Y�jf>ΧN�3���X����:.	�eP+K/��u�#/R=ۻ�=�<fd1��:E�y�����=F�����=��cP`�DkRj���Tjě�d�5��F�	���nj������
��E�XD5���_���eI�G��6̳l������L�S��@�tb���j���p֑���5�wj5���#�@w�G� Tq�pƉ0 ��C�y{H�����H]`����'��^㇨�w�㾤.�7*CJEu�k�!�w����>`���y��P��e���Fd�Go��G\F�E�"�z�
{�Wm�D��q�ϻ��L�4�O���.m�ͥ3�k	��v �m7};�.3a�0�	�c͓��35����������o���Xj��vF�r��B$F6�&&�ucMa�>��@�#�����t�G;�dMݜ]��3�P�T��v��(��� ��PA�7Ӂ����{��J��3����j����v�/���)�ߩV�3�����*�����u]F΄tT��māeVނ���f��\]����b���mq��LIbRȠTA��!��4$v�)�n؍8�2"�ְIFz�7������]p��v
�$9��g�������uvݸ�㣎����6a�{���<�:ⱈ����O`���r�\uX(��c��p����"�:�l�m>�n9�հ�t�糚���c���Y]��_Z������l��7ݰ��ۛ��q�	���H\ݸP/d�<w6��[�-�t����k�v�F{������*6J1�cjCQIX�h�m�1��PF�6�5����Q��(*��p���U�KTc�G�]ק�7\N��Žu��̅qƽM����.����s��>�3�
fN��͟��0��>|��2|�_� �����CT��t�?���	8e&nn����p����wgV����Y����0�Pt��� �AL�$F�i�5�ήtfJ簌����G���g2�ޟmU7zΰ��L�Q8�f�P}�D_�l���鼅�����Q�WOg��<��@q(Ì��en͇�����< f�UC���ܜ�_V���{Q���U��/��kvU�����;'&���벷�l��{wo�Crԓ�*�v�H�)�
)@��O���y���V<����U���>�V����Okm2"Nd����������H��!�|��B���48�p\���s'&�t`=`f��Q���T��hN���c�ꨀ�(��1d��V@�S�//y��7��뗗w\�r���P�Ѣ�m�,�
-IT��,j)� M��ٹ�s[�EH��[Y��SZ֧|�I���+*��x�r���p�Iֽ���+2d<�n�@� \�����gv�MCZzl׺oG��㐳Ê��f�o$��}�+2ٖ}��F�L�c�*[)��F3�k�b��i��⯩BP.SH�j�гXk,����L�i�>�ww6�a�w�䄬40�#�]�Mi���@ut.�C{�j�q£E�7��l�����vl=q6�#�S��j�<kk�a����o���K�7mY�S8ø�ʖ�fҙ�y���Ri����b���2N&��[1�u(�-�e"�A2Y�T�3��P֑s�|��}$d'���m,�e�e3���i��2���M'�F@-�Kf9���:�&Z*B�)�����ak�9��=!G�L���A�{@JѯLy���1�PP���9=}�
�����ll�F׊�/
�Xˢ�<�Bg��>���+n�쨿e#Rb����:�tb<�b;���[/�������#1��kz�&����r�p.�w7��~yT\\�.�|8F�=Z�wW���Ni�e���c�������!s��of����<��F;��3��۰@��u�	I�LoI�Mib0z�n��x�{)���}��<	�|{&�W��O�]]�f{��s�E�[������ȏ{��C_x���.���k�j��
��8���{�����-������1�}�FlU�jR=rJ������n�L¥����~�����Lpp2�VaOT�W>33nC#�#w�Ւ}������(����d[r* �g2$�n1����vF���-��F9�W�LUs笀��i�s�6��܋�CNu�Q�2wl��Z�	�z�ilL��>�q��XR�r�w�>w��vU��Fx,����N�~�퍪����_���b#���kt;ݑ�{y�w�~��s�	�v�3�/M�'W�{I�V:�Y�}Blٽ��3��퉞����㜕�@A��w�Lع<M4{ӽnx��L��/I��=���^o�	��/��_d�A$�=��o�^|6�mF 7��������Ľ;�_)���޵��{����_zO�qH��c<�2R�
d��˘s��_f�ya�|�S�`ݾ��it�r����`��9��;�_y��{�O��-���yUK(�KO7f�L�Q!3�8�wG�4l��]�o�x���v�:#�m��ל׫z�,p͞��Ip������R��ה �A��tM�0�)���E�L�xx�j)������/����>�O@�ϟ�����W4ڻ&NY�.L	�x�X.4��e�|���zl�����;��ϰz@���1��&?/����ߚ}��[5�f5�V����l�E�e'C-��{��5<���q�oL�]��w(^�K�=)Ś�ƭF��5NQ�U�k E�9^B7g4��n^�����f��%
n��'�>�嶬���r��X;Q�O�=s|2V(�[���夌��h��qB-���Ht`:p]�|tK\`OEC��{��qh���|����^��V=�&s�=О4��^�"
<�&n8�����g� Psk�D�Γ8�����cr��Z(�7�}�vM�=�o�S�Ǯ=}��������<�vO?a���p����#i�UpIdn��H���C*�nmЙ����ݧ��|S7q0���1 i[�)QJ/O��"�c��;��S�3��k���<�(F��bDJX�i��ur=�}CQ����h/s���Vtc���*�;�=l0뗜��D�ژ�:m�9�s�q瑻��^^����Bd����i%syC�����)$��$�=�3���cf��KN��]e-O�*�+:�T
`��ȫ�"E�Q���mr���ksTj��F��QBdU�<BM!I������"��z�@�4�#��Оa):3��2�L�~ `!-�^h�)4�'��R����S=�(��M� BRg��+l-�fY޽|j�i�9�e\��m�Ͱ���i��/�Hw�<D�5���l�l�g܃Y�4:(}��~F���'%���#E�+�]s�:������1�����h��w��1�|ss۶T��*�MCA��z0J�C29�0�٦e���t��f��w7��Mk�����$��m�L�*�M4��n�Y��I)�e��u֍2�U�>�̙u�0J�]����|kX8��O�F��&��ikMCK�ʃY�2��j��Ͳ�����w���>fѦ�����a�i}c���d
g9��e�l�-�} HZv��SiHi)��Ɗ4�&�I�s�n�i�m3�\{�/�s�ݯ$��)ְ+�7�m.�����*�#{`�e\anPטIȟ$/Fƕ��.�ޥ� �r�\.��_5_wf��5��`),
(u�nQ�kc�E�o�lkx�sX�B,<Hg]ԣL�����>��(T(����H�"�v���l���ם4L�iHs-��L�i���5(�e�Y�㳸^��Xˍ�wW�Z:��ޱɢm�Mn�6�k-֞�Kdf���6��K.����~�G~�s���i4�,�;�F�l�)>����<HÌ�q-���ʛg9����ǯ<�%)�
)@��٭!��P��0� CL�->�ە4�f���M��)6�m3��O�|G�(�5�5�O|�m�	Ǝi�f�l�)=�W�\�)�Jg�uܣhm� ��ZwG�L�IH}����VF!x�2�p!�3I��dt���z�z�!I�Rc�}�����1��Q�Zi��Ӆk�Ґ�CO�X���0Z0���#MNX�b撙�����a�2�g�L��,�+��6�M��������}��\M���7���}T�ca��s�0���U�ю���}�4������m{g��emH{�� ��\fC�&:Ze(C�E�#dI	���XV�wg�z���lY2���/��;=�vp@���/V�R�t�&�� �V�2��x�E3Ց6+�<l�ۧ��5�^�8A�;�"��sm�J]��4��l]];rۋ0Uq�^��L skv���93��̓Wq�'��<�������n�0�	���[>{v^�Y�����oR\�c��	g��s�����wv:667�r�ci+����6����ĄKlj5IZ+t�J�r�F��?{�n�]cU���ˍ�ú�>7mT��D����c����7�$�����qp7�����ikMCK��*5f��#C�54�f��s�w(�$�'��-;ez����MY��R�@e5�J!CcM[6�N纕4��ٴ�w���Ͳ�l�ǎ��ͦ��S1��Q�x �e���&H�1
Tl�i�kH����m�M��맭�O@m-|k�����u*ȄS5�}-�\fQe��M�,�M� JL��d�i2�9�i��I��RҒt%3}��$�2��Z�O����f�3Xi�_�2٤< ϳ��M2�e���v\����9ن���Lת���l����i��-[e�-��M���\�	g��n�{�����ݫ���6a�p�"��-��>5f�481^j[)�Y�s�r��m�O��VЃB�P��w�-f�<��T������e������d���V�~<�t����cX�H۸&~<DvB3l���p3�_1��EҡTG,���l�EmGV]Ɖ ��dH��U7.�����Fߺ��u������"�)"� ��]�oݮTm�r�����-��6�ŌQQ4H*���k����mw�����dz� R�4,�=��MDJP4�%����44�#�Dh3Vi�Z9�e��`m���R��L3�>u�[�ӓ���~�0�6`(7���W�b���W-�WZ��a�o~u*i���)>��׈���!}c�>���Tm��M�e�l��?jQ����������2ӌ�ǎ��ͦ��S>�ڔi��5�P�OJ_ QЋ1��e��f�h��6��}��׵�k�n��Ի�Il߮�1�!RF$\q��7\5p�kߟ�%i�#MB}�;Xf���S1��h�m�f�i�̩Xj�!����19"nH���!��Zm����kl��Fgl�{�F�L�)8f���)�Jg=���gI�&
��j�燯�H	bZ5�CZ�f:_�4�f�I��R��Ig2b�����]()rf����׻�M�+=sL~�Q��9����I%�w���%/n�8e�fϜ�ހ"��b�6��(���l�^���XȢ�����Rsp�j* �Œ�6����Q�1 ��X�L�Y|������e���ZF�P�y;�$�p�#f0MT�l�m���56��g�WwIsl��س�ưS4��l�ƺѶ[4�G<s�N�0Ha	�.��5�C\�:�sl��)���頻�i�e3��e3L�ٛ���S��<s���2��u^�x�]��u�u֌d˝��#�I���]G:�H��.��;}�o�����������I����4��2���F�l�)9��QЈm�ͥ���[�e��I]�^0!�7vkH�Zj��J4�#-�e��M2���s���.m��e'ٳՆi< �Ͳ��wAj �%����֚�u�L�5g9�_76�I��Ǐz���I�}���CXh���
q�!�:��gh[/���R}�Zm��͞�3IL�+/�V}�ySX�γ-�[d���s�סk�{��W��f��i�d8էba�i��v2c��.�����nb\�i�@P-kX�3�>�1������'UQAb���Ql��\4�
���ͣeݷ�*��-DEB"���ww�֩4��n�� K���i��4��P����5�c6�|�'׿%e3�������S4D5�Ol"�MYj�83ؓ�IRvV�u�K\U���lv�#���i���V�ζ��f�e]��aD�j�l;F�"��f:_�4�f�I����L�S=�V���)6�Lx�kl�i�e3���B�8�-�#"ƚ���#��L�>!l�[9�w��6�M����Նi)�e3/�3�	�m�şcx3FD!i�u���4=�a�u������{[f���2��װQ�S4�O��YXj�!{	�&�%FSn\q9��Vw�C��<�����H�/�&d�_ٓ9@^�tb�o�����db2����o��@ݿUS�	ޝ���<�Cv�qA�4龅���moFQ��]�(M©,�V�J�/PDz���L�EMZ��V��h�*��U��wS�d���hf����z����ٕ�c����"4
l��իX�wZ��m�����<�G�@��`��q��.�-k�l7��gc�Y�M��s����wc��V��x��pF�"u�#fE���p@Y��T@�k�m�g[��q�ڶ�<gǷA�\�:��s֎��o����x�>�f��d{q v�v�����B��:�˥z�;c[ft��.�^��z�&]ک�S�d����na�%d���d��M3EI��j*4F�I\HP�X9���PI6�۷g�WCŸ�;n��$�=�+v�����j,GY�?����P�"��bC�6yX�L�i)�}��b�ٔ�)1�u�m? ��l�-�_�fY�Rr���VW&j(��8��MCZD5�&z!u��(����4z��Rc��Ѧ[4�Nf�54�B�Y�4'z�R�F�r�u�����{�4�L�7_^
��	4�N|W�s��m�����\�-�S};ݦS8��1��9��m���L�K�P�[2�g��e3L=��n.i��`	)=�{5�|hi�k��ƒ���Q��q�t�4ӟ��2�%>�0�o��.q��e's~if���S1��h�-�e=�=]���7+�ma눵Ĕ]؁�Ӹ�p��q�7u�Y��󏯱��<]Dra����}��{5�G_z��0֚����Q��)�e��+]nm�ͥ3���~
6b�@Y-ƅ֚�4�#���{�������w���S�b��3Ϊ&�6���q��F�v����
�F�?��ݰ�?ڴ�υ�=���1b��7��%wU����Θ���e ����L�A���Ld�h�ܝtDhwn���0�&4_�e�L��l�SL�i)�}������>I0ai}=���"�&PLBSwf���L�'�	A�L��s�)�ڠi�޾���5d�x�iq�.r-Db���Y�����)��C��m���'��sZf�< �Y��pP�!t��Jp6��6d�L���4�a�Ќ;�y��a�e����L�e9���S4�ϡ:|l�\�c�Ba�.�a��pp1Ņ�:��ĠCټ��>68��W:e��I�)2�r)!W_�|j�߽WL�i�e3���F��i�����g���-�Kg{N��6�M�|k�Û0VF	m�;6E����
�÷Ń�2d�s�V���;ٳ|*��a��q�d4�j!�vw�<wf�q��n�E�9��-u-��+"�?�1�yD�U�b���d��S�;v'�j͊�rM��kj@��<������s��W��1᧌��z_8�%ُ�kz7�P&�$�E%ň�v��#A0���"���	 �EZ�92E�<\�ݳ�@p0�B�9�Jw���H���߶��I�R{7���M3l�s���L�4� KNv����P֑w��8�*4�P����)>����Jf�O�g�{�6�f�I�l���S4��������I�B:���]%)����J
���Ǭ�;�����pՇ��sZ�[[����}�L7uM�K��#|j�ύ�e3l��k]nm�ͥ3����x�I0p֑�XG���a�iN&z#."፴�lHli�5��v8ea�P�ͥ���t���I�Rc��z�M3l�s����g��q��j�����p�3$l�!��P֑{��j�MY�!w�	�"� "�՚_�k'-�ɒw�q%�6�('![�{B��g��}�'>�Wc�Fs��c� }yw�6o\�;Ȋy�^\��;ȚȾ�ӲTʗ�� �{x�3�\*+�w�nKІ��k[
~ޱs�މ��%��;XΈ���oX�}�ɶa��X���UFD;�",F2wn�������a��Թ�Zm�����!�'!#.&���/���̞����ϧ�ݴ�f���ݛ�'�������"�3s��`XX��7����7kg[-�l\3wiBw~���mj]3�h1���ʾn���]ͽ/��1sjK��N��ºH(�!C!��$�v�u������+��Ҫ���GWo�U��@|/���|�l8XP��V���4)�e�i�ވ�E��.�>����[]��,!�5�o| B�����ݞ��ٳ���[��P_fx�ْ��.�"Z�CE�i�5��s,�ZfY����L��x��̤������i-�e3V��6�f�I�>����^N��L�r�g�1O\�	F6��U���b���W�m���k��x��K��=[�kP�	[A�.6���Zo���Fu���=	�Yݗ�G9ɘNc�A1g����R���H��+0��CYnf�&�v6[�;q��1l'6����׉�H�:�,��y;Uя(��q�̟-��]�mM��L���vm���eY�f�"��IT�LD����6�y�ħ{�;@��Wg,y��X�ja{���Ğ����7fjW=���9�\8T8�x�p�Nw��V�3��1��r���-It����[s\�.�
��S��k`�H�|]vΎ���4�j�R��ݻQ'��H�ᡲ��ޗ��z��8Ϻ�#�%�i[]}4'�c"r��LQ��f8��W��W7s��>���!LV�w�@\��ǁٶ&
��Z	S�dn������[&8Ƭ��b�·$^�B�ݔ����[fi\�˚������F�ͽo=�~y��h���!N� Le�:7�4�����b�栉��Y�,!�=G�'lg6��M�$a��B3J�n^И�v��h-��c�'�j�7o@�[L�7\ĳ��g/�qp(.�$°F�X�N�(��}�� :nc2pψ6MԔ���l=۵s���# �		�#6�t��rf�#��"��!��W�K��#�L������(�:s鏱�����<��>>ں��%
C�f�MK����sۂ�KV��[��*%�p]UT�obj�nHa����`����S����1��Vd�W�)��F`�a��S��˺�Y͎sZCn�Y<�{<2'��ܗC��|g�3�g��y˓��rhV�k�r�8���%m�ۆ7d.�Z����W\�9sZ�wGm��]��.�%�zŴ�0*���ƻnw��$l���z��Yw�;$)��]�t����.|�]���m�k\v���ɧ��[j��l�/m�@ul�5<���>���l^(�ǵ6y�x�[�=�����b	A ǜS)�΁�.�=�W����p9��ڕ01sC�m`�f[���6^�[�]m#Pn����e��wus�M��A�%���X�x�sL:.�ƻz��ݢy�n�dˋۓٹ�n�k���>���[�S`1�2�8Z�76�;g<�9���Mo3���vA���5k\��Q�./<J�{nM�;.��n���p񳂻�ۮ�u-�!�׃�����96���v�&z���ǳ8������G��@���:Ćz�Y9Su�fǣ��<��t��mh�:Ѷ�b]�nۛ;i�1[���2㱱B+���[ll��!�q�rai�OfNګ�rs{<.����E[�{W�%�c�R��=]�v��p��Ys;�����M��vl���80޲u��A֙s�B]Q�V�W9��n<q��}m�\;s�lQ���^g��g����;��v��m��t�mҘݸ�i�wM�{lv���Jۨ��E�T�Z7'Weؔ����P��9,Sr���a������!��].����uƶ��U���l�=����pq�Jנ���wgzf�f���i���tu.s
۝�]�+�q<�K����j)�(�ݵ��ø*9�c�]3텭�E��՝����Z�[��*p��]m���܃�n�z{d�':k��+�V7Oc�����8Ϯ:���:v�z��[]���j����mWU����&�{���;�5�Nc�8��t�uǑ��k��w4Z-�>�Ȁ��(���K�����9�p՚��\�U�]���zlquźNK�Y:xv�ٽ��
����Pp�`�q������-�}�pǲ%�6��C8�� `<���{�&&._^e�گ�&E�͝%��y����΍-Qv���š=f���S��<��z�iF�w46A��j.ӹ�����Y9�{��3f60�n�B�a�0��>z���;Zv�=�u3WcFl�wnʙ�����r��튁����Xa�Vٮ���@�@q\0��ڟ�V������Gn_n.s�;�S���;Lً=�au�g����+
g�mMo�^3�l��|^>{p�EW��!�o6o�������e|�ۢÔ��k�Kk�wZ�UW�x���-�zP�=��]�׹v�8��-څ�0��5�U©�Jce�:@)�9�\�fS�N@����^�y��4ψݺ�-*^�K�ReH��<���ﾨcEf�pw3�8`���@��5�3W�K�{�i���.����^(E���'�Q�B�h��V���&ɭ��R��+ �t
3D��`�#���n�ɡ���^ш�&�w3|_˸��6Yޝ=2���LDg�sA���'v���儌o˱����R�Ş�
�k����Hl¾�x9� ��ډ
�b;� E�7<7���f��-�0�2�a����f�����X �ظ�t��Ð+_�(JFT*lK�)h'}*ň.���L�L��{�aj�~��<�i�X8��0��"��nkϻb�g�qv�� �qtvø��<���V�s�N�|]ѣmǝ�b�;�A�Gĩ�c�[�o<m�K+�۵\���t�a�ճهcq��J8�X���)�z�n9��˻���>��XZ�6�-�a�5x�v3v��n�W �`=[g��&#z�v�vݞ��vh�+ssۆ]���ZҺmvܯf�11ʉ�Xv�Y��p{�?gn;���N����Pi7wd(/}���읷᷎zp��L�&��[��w=�=�x���-�`{�2c��$7Xj�!�>�]i�#MB8�,�L�)����=-�o3,�->��L5a���X>��l�"�u��e&=}�e�|f��[>���fٖm���k�Ͳ���}���\�<@�2ӯ�}p!J3m�&��kMB>7;�Ѷ[6�O���SI_H`�[=��N.q�v_���a�5v���
���#�b�^ٖm�"�z���L�S;���sl��)>����Jf��[/���6�f�I���9YS5N1T\�)�J}�wN,�)6�| ����]3��q���sz�6�Nv����L�S=������vn�����I90�i�n`��$ۆ�h�V�.۶� �S���h�3�P��k-8�N2���4�IL�S+�}�4�M2���:A6�ͥ����V4�#MB��-�S�DSF�}b(z�1�ޛ�ŏ��Ȣ~m�Q���g�U��Eʚ�Iq�5��ݚ8 Ǚ��y�:Y��"�5�(]�N6��a828�J���PoT�_+��U&�{����}M��h����q��,UbہX�șaI�޼���Y�ױ��I�e>��ji= Kf����(�r4�1#������z試L���1g��D8�L{^ǳa��6��{^�f�I������eqLH��H�!��!¨����|,|Eje�k�D�-2�8W�i�M3��>��c�3O��zQP�ӒF�M��S#�Ǿ�;a��6���׷,�)&S�{<n����ru`�DxUw��a�E�7c��Н�����+��]��Y�]b9�̽���(șąݑ"��BFd)��+�3�-�@�8�R�0�r��Ş d�L���z�Y�"���2�r9�FR4�@����4�H��;��,��fS�������+�}�4���B��;��Y��
RAE��"4�k���V4��P��W\H�8�g~�g9�z���}~W���Q�$��Z�Y�3��$�Y"��}z/.����?����v���lS�w���]��&2�vN���pfKw�ƌ�~cw{{�?hIID��4�I""��	�;���e&Ф�k]nl�@�!������,(KN8,i���OW�(6��%!_�ѦRi
Nr�����4��N�z���-8�"ty{
D��0�ƣ�4�5�D;���e&ЧČ�o~nq)%3���\�-6�N�)f���S= ̾�k�;=��71�L��Hyܫ�:�z�]�5�N
�r�^�u�խO�[���k��i��l�q�Zw��%M����w���Ͳ�l����OB'��-��{rͲ��Q�ҁc�8�E�XrCu���"��;$��-=��K4�f�L���h�)�e'9Z�T�}�6��g]LO��n(��MB4�#���ikl�}�wrͲ�H'i�����)�a�=�.�՚�ߺbq�N8�-�&m�� bS+��5�ٔ���M2����w�n��!<	BA���ޏ��Q��3�U� ]6k/�KE�7ۂ`O;���,ȱc1JS���I�L�T�S�bB�t�b��乍���5Q�n��ǵ����lQ�j0W�tI,h�i2F4�0�;:�CZha�k��+�,��nB�8�Ըe�fS�W{sl�m�����6�a�����i��(r��5����W���jDK*�LIlA!P@���wsjM[���j^z���^�J�յ��ɉ�Ź23T�Xn|��}��Kf��N�q������sR�BRm
O�^�֑h{�ǭ4bQ�2�����!l2��u(4פ���Mw5�������e3L9�����v �
NY��[l��
I�J٭44�5���FY�e>�~��RzCN������e02=�`��i�Lj?q"��d���.f�����᩶S4ý�t�4�M����g,�i�OH��}K8j�P�\�/ѐT1"Sa"�7Zj��s��)Sl�m�� ����ͦY�S>.��4�f�I�V��4�f�������{*�Ɇ�/x�w{6W��{u-����``٤��Ox{�l�� �ZD�1�q��]�#W��gfҠ�%���Ԟ�}�	e��(�h!���a5qs��/�sn�4�;=]���/Ur�]&�����7c��;�1�wJ^ڮ����=%f�W`�4y=��R���6V�9��6�OA(��U��˸%W�ŵ�Z.u�ҳqC��{E�$ε��ě�ĺGaG�%͵�Vgף{u����\x�8ݶ�xλ[k�K�4�]wb5�M���3�.�Ϳ���q�$�N���"Q��H!�ܐc)z��~>`v�����h��JT�6`�-Y�e��gE�B�՘�V1=B�8-c���)6�O_q��I�i�Ϲ_nY�S6�G�����ޫ5�;���Og:=6G����ײ�w�
�E��VG95+CXD5�LFV�a�B��Fk�i�5����a��*%IIV4�3l���^nm)�3�wytٴ2���`�-;��m0�a�]s-��)���[��l�
$J�+9B�׹x� D�)1��1A��i)r�ܳl��; :��;����"��YK�"(\���͡��)=�{X��e�JM�|k�M�i�)>���4����߾��cMB4�#�(;=����F�%��lwC��p��mv*����mUӜ+�y^���zߟ|���*#A1�+���_w��V4�M�I�ֺ��RJg>�6i���Q�;s��m��,����%A��j��#��D�7{а�+��ى�Քz���ᅚ����q*+B]
������e���*o7NE�0��5�3�9ͽ˅w������T�����#;�ׯ��� Ѥ#�[���D�(LB0R��|R��}��6�&�I�_}��m4ͥ!����6�IN!i����B��Y��d��H��5��|4��M���W�A���6��ƺ��Y�i���+H�"��H@4�A���li��(Ր���v�a�JC��nY�Rm
N����ҙ���>цƚf�!����eDӎ$�y�Ͱ�e�+�M�I�S����T�S6��w��6m��e&=w7L�i�e5�3�������h6�����{n��g�Z۝b1-y���:����/��1�Q6܄5Q���k�P�zg�֚���k���u������@����T�XkB����l%R��GZj��{��e;�KN%�=��7L�i�e3��nY�S6�N����Ӟ�bi�&��?,p&TE��$.n��#MB:�z#XD5������®E�9�f�r��6����[��qSR�-|i?Wcס�Y�h��똋˻���M�s��\�����d��4��i�bz��5Г�u�)�L�^ˠBRR�1)���ބo9"*];�b���A:I��	((�=��o���5�����y�������u��|/��l���H��F�*�k4՚�9Ɉ�ɓ����|9�e8�Lz���3i�m�Ͼ��ox�ꯈ��#���e3D(c6[2�,up�>+g�t��n����ٛ<sj�~/���Ƌ
PHI������jޗF�6nF�Y���ǈ�ɒ.u��[$1�Tװ�s�f�P߮��}[���y�6}��wG�xЫ�vǦ��r�0"��l����Ӫy�W��DD\��#1[>�[��9�;��M��Q����P�M���ox}q7fޗF�U�e-����;2���2Vᣚ;,�!�^�æ��gݻ��Kst�C�	L'[#$���,Ys�:��7���5А*��-ܼ���b�^.����{f�`�,PU>L�����\Bi7�Ƀ@�(�585d̚;�ÄG�&AAz����wj�����X���wo���L��
�!�Q�RA���.2��n�Vnzv�J9�7-�is����<���<� ��1���_:l��4��g)ԣ�`�ZKg{��Y�2�e'����M(����E��a�"9���f�I+��u榒��S9�ݚl�M��پ�����Z�ؾ���F�`�"���� B;�r�a������f���#�Zc��=t�&�c�w}qB�['�p��j,��t��!���_rT�8�e'�~�3IL�)���b�2٤�A���ܩ�S4��;]A���-�1!��L�5^���3n��O��w�m�fY�R}��SL�5�qmJ�ZF��}Ӿ��N��݊U�P�? 6T��/�^_c�([�ښ�c )N@�v��*�/^*��h�o_D���̑����F���]�2�U���2'M_�Q���DD(I�pi��v�N���7嵻[V��L�&��AmE��C��좋*n���D1�7p7h��^\�Y�"3�]��r�v�ᢻ	'6���u��\�F��<����Y�.��{.g��m��xx�^Ύ��T���T6�mk���	�֭�au��=op:��rrb�{i�%$���:�c�Xi�>^Q�up�����9�H�NI@D��of�bJ�{��^Nyz��>��Z��kn��=�d��8ۥ�v�ӴGٰ��rkS�ĔvVm���{�tͲ����(�-�e'3�J�JCIL���g�y���4�����٤�;dΔ����!��l�cM24��4�hm-����hm6�Og�(4��%!���(�:��i��}��M�"R��%]i�f��鱤V�i�����i���-���鳌�6�G���P�r��8!@�*S�<T��i6��-=^�N�S4�f+㸣L�i���5(�Z��;ޜ�s��m��:R	�[�� Á8\�kH�Zj���ͳ,�)��Z�Sl�m)���ܩ�m6�Og�)f����<I�����{Sn ���u�r���zvqu�DUJ�8�8w;�W�l�k\0�;��-8�w��Y����w���Y��L����פ��6��{�:�l�m'՟.3�#"Ta"�7XD"���n��9��t�n�i|8f�/p!C3��Uּ�X��͸E�WH���ЂtS�zD���M�Tp1
^E�1li;K�-��������wLt�t�c���@�3  �3Edi$�eHQ��1Q�F������[Ĵ��Q�Zi'9��KO�/�W�K��"�B�%Hb��V�d/O/\0�i�g�}�Vm�| �e���Z�e3��}YR�Ց���������&B�m)��Kfo��F�l�)>��J�e3IL��m�.m�M�@�ZW���ѯ��Zj�>��*&�FF�Nlk2Ͳ�����e3IO��w�6�t햞�vRͥ3L�b�=�4�M!I������T)�G(�%D� W(��[����\��8܇��<�[�Pn�Ժ������RJg��śC)�Rc��w6M3iH}����fi>�{�JI{��W��6�P�N�i��}���i�JC|v�2�I>�-ʖ�`�w��]i��D|j���EQ�#!2��*酳L�;ޞ�l�6Ø����X�fe���}5��+�#ԉ��OG�ޫ��sald��-<�� ˼3l��l>��{�Ξ/��y���2�D@P��l	v�M������=��e��t��N�<O!�%�ݛ%bw{�!w���r�o��ž>�L��ߠ����ȁ�/�\�/���Q��wr�u��p�O��X�O,��`\��� Ȧ�f�R+���o@�X�+�%�������nw��b�W�Ȗ(3S>ʘdl⍭��c�U�ΎƢjJ�]�]&L�(f���s�B�jyvr��:/��4G9�K2d��C*]��b#�0\�܋p#0�Ti(�sc�0y� ���y���'��a�A�f��.>��ڧM���[�ޜZ�r;�d5lG��������2-7�c���/�ؼq�b��y13v��ѵ����P�^�0x��`������¨3�'���{�׹���i{�GuI��nD%�32F�+z�i�0N���e�td��e����6�-�~w�t`z���=m�[_�����"t׷:�֡�X�N����/+M	�ܡ�'&2VЅv���u	��呜o�����yƹGNfT+j������	d{,����_=t^���:�Iv�����%ǃ]�y�˥��Cgf��o�)j^ޖx�V_[�]��n��Wp�^���m7޺K�ｃ�Wc`�b)VN互gfTf�x �E9�*'�9أDy��L8�^W�XӉ;rUV��q����µSɽ�d�o`���Z��fU�ګ�������r�"��S�_�ž�7Z�N���ٴA��A������9+5�	�DiU"��������)������N5��ը-��c�ݻw�]jME��`�i/NS:�Q�D�U�(�\]y��z��ql��83�-C��`���b������Tw]���f����Ót`h?5tƱa݈B`'&���<1%}J�h�U�K��x�i�pL{̏�Z�e<L�3�7���۸�t���`XrQ�Lޝ�4� ;ul=��I�7���� Ѳ��Mx���FM�L�����׻*@|M�2��2*�{��;��~���{��g��ٷ�܃"D}��³b0VL-����#}�i�9����uBk.[��a�'�:�h�wrnT����:�V��M�:��ԁ�����,݄B���m�PYJix��3u`��e�Օ�"I	�5J���-|[2���%�^�qlo6���N��N�x�1��*҉>�	�G<���3iڄ/n�>�5��<wq��mE���{�P��ǜ'|�����1��r��pw
 q�2;�s�z��VLZ�b�Fi�xcov��<
'C���@��8s3� E0�8ʭ��^�Õ�tU)��ϧdX�Di��
�����������������w�����O{��xf�9����t�B�	ݑ>�`-��^����*�z�>���g�s����F�NQ�n�_�ۺTI��s�QF/~��nd�""�*�����عSL4̦�����-�g��]v��C���g.\���q���J�e0�;��{��a�e1��;t�٤�L�zz�3��-1��s�ϓ(����u��֑|���a�#C�G���Y��m��WǱF�l�\�:�ɓ�P��{�����c��7$p�qV�.H�띔N6suù{v��sݭ���
A��L��|i��B��z�#k)���⍳l�)9�뭏�c��8��_q�,�#M�|��"�1��Q�c8̰�S6��+��F��&�l��ܩ��4�ϽݺśC)�Rc��w6G�V��� _h�x�TI��5p�cl���g��sihm)��u��H[�A�->κ�Jf���|{i��AS�|�i��J2�u�B��-����b�!I�Rc��{6M3iHFxX�P�#=�a\��p�8V-������������yH:�޽'fgc/���3�w���#�t'�aX?-���w�x���7�+�
�A��Qb, �ʍI��a5�鈍�A���=Iw��sil�S>�8���l�!FB��ȱ���5㾑+���-�3�e�l���u*i��}�n%u��j� ?b���TgX��z��f�gK��^�z��rgN �5Jg�����6粣D<ݬ�'�g|{�D�Kj�P�{�oc����p���!�#��a5��f��y$-�Pa��a�G>��V�,�F���{�����#���FZ�Pֻ0aV�Ց�O$�T$FH�9!��[6�ϳ�jQ�Zi�����4���;Kf/�أl��)>��J�Jf��Y�_:�q8ʈ��ƚ�i�Ud;�qSil�S9�:ѦRi���5���ٽ�E_'���tvaq% (	p���,�d̞�9����a|�nkt��6��iá�%��+>��*��U>&�j�Uo�zb���!�ը���u�H-��U�:6��*���SVmE��V���5�#�^���@%PwGqq� �n��7V��)c�>"^4�gÂbv���x��荓Zӻy�z=��5�tuӥqj��L砧��8ɻm�م�V���P=b{=�ݹ�ݸ,gc/M�v��xu�n5�GcSc�n;F<�%��q�v앶V⣌#�u�.�;\�U�9��l�d����FASk�̓vsn˺M�7R���5w)���bN�N��^�u\>���^���C$QI`���	�v�l�ۙ �N�I-�  q��u�>on�5���;6k�r&�f8�:˷IG���s�ۮ�j:y䩜��
�T��_[���xxת�����ۓyg�3��.%"jH�I��/�lu�ޱ謇��:�o���UO֍�
G�����W��6�QN�ogb�ЧM����DD]���K�ڶ..�rz|�qD�i�LH��n|*���x��|쾕��ypf^z��o�fFߺy��\p�R��ݣ�ŵޏn<��y��UV���F<�����	`�F<8F\e��tZι,��r&K��m���j9x4JPS0Z��cc��UM<�f3H���@m������;g�08���� ��n�}�[�ߩv
��pM�^(�%|������G,������䜹ض*�mH-]T2{��i�J��|���7��4ڷi�9��	�D$J�1�ԚK}6�J�h$H�%�d�A_=�b�I�翓�)U;�Z.ݼ?�W�芹g�y����$��od]��2��� �qldf;aw}n��}���RI�Kl�{��W�M��鳋�+2�}8p�gj��|��2�8�m2C�d&Jݛ=�ѣvl� ,;�}s��N;��'�yïvt
}��a.Qm�b `H�u$4��6.{O�h��WŨ災�Ѻ�gn��",�k����+ٓ���UM����S7>����_x�4n͆t�3��m�a)@�Q8����<"��z��;�j���ת���U�4�Į݃�<��(�-�	2��v�J�y�"���k�n�WPn�d\Zp;�j��'��D��_�[8�g����(�W`���ѐ*&�֮�c3uU�t���|�};�{[/��|��8�66�э���h��"eIS1h�VɓA��
-%�r�b�߭�S�շ�tE*�����Z�ڒC�w��mn�N+�̙"�ϖLΈ����U-�(A�CH�.U�c������93�kݜWÙ2j��̼��������\r��5���5��:�(�=:ԯY��Qt���ݨ�Ѻ@l8��>4ꝑ>�r��b��z3'$w}w��wБ�8[���a׻9ם;�U��|G�Y���wL�MY� ^��g��7q�#L�]n͞��ѻ6�wf窀��<F�����׻=�1����e�c��� 'y�;���v���DU_�|mu�?8�̏�9R�j�3����ڜ�{��F�)�o5ݍ�)h��]�W�L!%�5ӻ�d��hw_e��Y�m>9����8{�}��,YQ`�·H��BTEPh�64�{9RXM�<sE�`�E��̦E *��歳^����v�E4�����ݥ���3�z3_u�������Ù��
�%�z��"H)��q����9��3m��ݑ���l�Ş�izz�&�6
l"R�J�v��T�wP��j�����{1�O�e�yA\�Y�B(4���O�~�DSݞ�T���T��C#4�>υ����L
	�v�Ͻ��Ԋ��.�n��:}3(��t�n)�JHX��z[Rr��R�n��vohj��?�͒z��'єڕJFF�����׻<(3����}#2d�c�T����Q�kv�՘f�@�[���m��JB�5#f���S9�44�Û����,'��ޛ�)�#+s��We�7X�Ȭ�X]�y��@6�^�M;� &A����MLz������h��J��6��`��te���k��8��7Mͻbَ��<�N��獝���9*����K�=��*��m���y��y�&��.���{d6z8󁥺h��έ���jm�vxgv�ӭc�m흷>mm���.������C�ZN�t�ggm9z��uf��y�v�;�H���t�»s8�Lg8�b�����Q�)-�ET�Ib��[Dh���h����b��F������?���2�[.���GqΈ���F�:���S�n�۬�EqV�F��ۛ��~����b���w��[{��G��cϯ���vzǽnB])L��R�n���}�����V�N�vEWG��N�y����"(
'>�����B�y�����FV����i�|(S�ˁ���*Cp(a��� �a�ݙ;ލ���yN�l��P�w�������߈��"�
5$�vl��f^O ��ٲ)��ə>����� �-at�S ����-�6��B�և<=�W槰�@�{C�J��+���N&*#jT��.{�w-n���f�p�=�������gq��/0a�b�yJ����>PGV����N��v��	��qs\���,&Nh�x*�$�D�t^efD�rg}ò���͵�x�]L�����f�s�Wl�����KF�71h���`ɬj"�b��ZT�����%Q��"�X
+뾷.��WO��c������}�${�Gp�\h��8���*�??�K�$nG���Q��6XR4(����}[�~Oޙ/�':u����g��z�R�1��f@[��ݯ�?�ITDA[Ѷ��H�J��9wu��:��ҐH5"�F܄�pm¯^���G��0۰#oP��W-bKD��V֥*M¹���|-]�}Ɲ,�1���E��|"d���W7���D�3]�:'��:��j���*������2#���O������4�f��T�艜�N.����|����6;^ȹv��F��Y��b��V�<�24^��&�c2+���ۛ�z�Ry�S���$E�L����Y7�Z��AAb��b0�b��wF��c�Z+F0\ۆ$�DX�b�TW�ś��������\j�b8i�
�ފ��}��>|�U��Fh��Tl���2�pI�I(��cz=v��W�𙡙�𞊮�����NB�H�P �A(e��9n�\��Cu�9��]��nb�gP����n���Y���c�3φπ2E�����~/�&�(9FB��fG���ft
����������z#��1�|�04SBF��$�;���lݶ�6�j�E��.Z׼U p}���~�.)Ӛ舱��ft<�U+��p���u-��M��D��j�押RwB�?@�:���;յRDq��4��0�� {	�ɷ()Z�4S�vp�
�A���f��V��a8r�g�(B��E�ɯ�{�"!#ҺQb��ͷ/;��h��ƍx�-ͮj���I�Ƥ5��lt>L��0[H�ᢜ�Ww�h��{޽�ww�rM^	��D^рg��\l,뛥�9����'O���������8X�l=��١r�מc�[���~�~~|j?ݭ+��)���G���t�2�� ��E�S@�w~_{�4�e�Y�Y��1���#���>��^`�@ŅI�:�Va�"e�����e ��\��0O:$p�"AȊh��UEO��=�f8}v������m��c���dh2SDfG�_:V�U �{�sif�&f��5R���E�Dem>��j��s�c�d� v;�����W<�B^�$������F���n����Fn��쇗�n�RY�_c^V���G�����e:��z�R��#$��*��X���� ��\���'f�Vl.Η�����p�]-ya�*�a;WA�x��U�Êl��<
�pxS�#w=���I�^�r��a�0��Pċv
ѷYz�{;L�OGI ܱJ$_r�p]e����$�5�nx�T�7�,��qN'&��d���[�g�^��{�5z'Z~������*��gbs�ڨ���`�Zc���)��45��޶�,Rr+5���x����a�!ǎ���B��G{w�GpMԧ��>��N_����u���5w��g���tw	7��Tg��%����+=\g*���W;�~��D�;u�!l�I�De��7�����j�j�^I$e��_���:p��uWؕR�c�r����pA����YL\T�n��'�`0g���{�C`�lW�c
�VLw�i�m������[ݼ��yS��O>y���d��;��ݻ���1���v�[�|(M`�Wf�4����9>��⎅u'Ni�j�aq39{��8�+n�b�z<���CK���p?kدv_r�&}7��[cp뜏����ݓfnt�!]�p�����1X�=sJ����ک��� ����њ#EmE��Hͼ��'���;�jf��oA~��$0�5��d2M��i},����'�j�Y:��s���L��5�N^jɒ�[�p�5)Q��uT�V_��~�����8�q^�&���:f͞wn����Ջq�gTz���. �G��(rpw��=pg����oDx3�c'pjk�Q��Ϣ�3�k�8�S���8�u�r�D'��}�ju�n���]I�ݟ����kp����1.콮�3������ld�]/(��>ْoC{Uu�,��+[y������oA�]z\�����њ�'�1��t�l���ӻx�w����w]�:��Ź��۰�U�6:U;s���	nnG���z�>�7���^��Tⵣjva�ဓ'\8��:2mizݘ���1хW���r��b���x��x��a�[vk��B��K͉Պ�y%6��\w=@��wGuy�Xy�nƝq�\c��Ύ{��^�g�����v��T�s��MVBS���ؼ)�4Og{G=wY��ι*�.2��Z����<\)�q̻=�ڼ�j�X��l�b����ַ[�ۧpi��z;n,qʻ=�S���)σkX֜�f��C0��z�Y���\���	�u��Z�|�v��/e�v�u,�c��qH��o.o�/m�G�p��k7>��nm�F1��W���tx�9'��x�zƓ玷7����������뱼mC�m��r�Y�i����tQ��N:��>�u�q���,w9�gu��L�6�����8vMXaٰ�����n�W[�9���6]���i�W�����u�vn�\pq��ӡ�wݍ<l͸�]e��j�q>-��n�ku�4���}i�n�f�64u��N7��k7�,�]��]����`q9;n��]�Q�S�P��wŠ�۶���.л]����u�3��-��7���L�ۧ��m�ض�Qݢ�-ǵ����6NF�������>�!m���l�Zcv��Gn*��qij�psY��ݮ63�F��X������pn#>�s��^8�ێ')g����敘�"RK�oBi=�x6b������sF��puð;Tyς�`�b�g-<���8vwZ՞�	��}a(3�\�����lvw�r5dM���$��#��>�,+Zg�[�;�iX�Y�C^뻹����6#>�8�7:ٸs���4YN�W=,�R.~��{h��!ȹrf&H��N��*�&��3K�12j�pL�I��w8H��#	����w+����gc�#�\�@�KLa���46Hp#".���3��w��:��ԍ���=%��%���Ep�{�n��,���	m��� ���K�AAyz>]�g�����D��Z��E]���芚L���q"Ż%)�"m��q#��cj�1�k�t�F�`F�s�psUl���z;��,|1|nn{���cz�ɬ���O%2y|���G�+<z�o$"�ӂ�u�0�c�K6!0Y1#ȓ�I��no��@���xf�s �4x��dQ�!�)5	i�rP׬έۦ����;��)������E�. ��_jZMJ� 0H&� iB@W�(cO�Ĳ�;r9����n��}�`�eƈNCGwE�Uj��è�����q<C��A*�,Í&��6�����݌]�2�q��c��qxp�F\��=|y�R∧xލ�q�SS����E{e
gv�:Q֮�l6�k֬�������X�$5x��\����Z�s�{`�^�JK'W��H.�.���}��޳P�5��x�o%S�ɞ�3o�o��h�o<�/7�0���{Ӿ�i�LS<-�9�=#�m��r�wWn�;�d�.���\j���q�5��]�K�6R���׎݇&�嵪ZL�n����vT�m�h�bvbL�0	�2��x3k��㣡�z�Ѧ݋Y4����⩶|<�mp��9CNM�u��ٻ��v;qN��ŉ׷\us����i�lK�7Z;WZ9Tu���F���ݼݝ�6�6�VMqۮn���z�v�����g.7Tq�g�᪸z��9��ث��zxsYɊ�S%%gi�ɑ�)* 2�a"��DcFI
�3����bݎ�px;��]�y;V1h���iEz㛌�x�BC�h�-�N�Iͮ"�.�8H2 �M�(�%Cm�+D�)��uY�H���U/�w��<�'�%�ʅ*M����
���\p�g4}�1��� �b��h�2e���Ff=���z#�����2�o��I��$ꄴ�Bb���p�������.��Lela�=���".�`�= �N	D$�4����է��=�]�k:{�ݬ�91�
�w���qE,0�Bl��h�k��v��:�;(��n{c���uf|��g��2�%��8A आc���\�̢"��ܾY^�[6{�[��y~�c�!i6�E	��v��p��'{"H+w�^�_��g����3�U�� d�LPK��
Y9�V2e\N��L]��8]`	�ީ��<�F��&��qb�ظ����{^�p�DѓE �ђ��s�DA ���kN���8rd�p|��(^���쑖�Q���gvo�?0j������ޏcߩ��+;��ݯ�w[��i�$�)	b���>���Ati�+3*���D>���!�>�C �O���m3wV����+�z#;��gψ��rޯ�s&>�?u4dcf���Y����+��=(*r=5����
���[E�Q�d�m��qa����ת�n��4����ވ�ɝ��E�����a,HBrC�{>F��(^_��X�M��|i�<�^���[��@�T �F9E7ݛ���sgݸE�Ɋ5��F�%��cx�]���l�ġ7}z't���(��ī���s|0��5e8�7q��Y�f�v:� Ǝ���u�;�R�y9v���S��*1I_}p�iFC��U�1q��`QFE���;���5jq��^`�@����s��s�����/�sE �=�m��'��8.0hQ��G�DF�L�9�q��뗀W���ID�8�NA�r\W:�m���%N[�zܵd3;t���13���R�PE����A��wS�J�d��{���t����!k���m��}v��|(W������[�PEU.�{;T���/ZR1bB'>���\1&UnV����1��MY�N���z��6H��i�{������= Ҥ3�뺳�g����Y�ow���7��f���\�ʉ}r^�S�q�j���ύfڪ㪦*�G:`)��*W�]��jdv�:]��4�<D H2�¢f$3FĐhѢG�.ȵo{iy���C��l]���k���f��v��>�uO2`Gd�PGSx)�$H�^Wぺ;nͷk�Sr@�8�M�X�e�;�j�.�Z`CN	D$�;�X���޺f������fVN�>�r��#J!��e�	�t����<(^��B9�'����f�����P~�紋�4ZiA
����gs�f�����@e���n̑x{2fE<~<p��	.�������������呋<*���������PB\-��q!.���s�2c�c��-ݨ"��l�J��ߗ�a���P�$��5�c�F\k)a����Y9�4Y��]�$n�Zr�#u���۾��5�(ؼ���I�k�(qA�ŷ��߭���әm�������f�e
�����]�o]�N�m;��%�
 gpvgZ�1���v;b�eڹ�3�,��4nN�=��7Ob�rݐ���3�ŵv�3�(7�����h� �N�9I�ԋs�ݱ��wN����ػ6��w��3;�얬����#��G��$��kO��Ƹ�ō�ǣ[���[$�鬙9����O��$ڍ���ـ����˘f��FF�����6N�q�n�'v-I��nf��8��]���/�>{s��3���+�M�X$�1*4� �
B����~L�T�g�U,�&?=�t��©�D@ߺl�S��eN���]舻}��*g�>��k�������S���$!Q"ѻ��!0Y��%tDEG�2�n�A��q��Ԡ&6��@�r�6����fU��O��ךj���w��T����Au
�\;�Y�n�UP�9���N�J��s/;@G޸d�(�5�[���zl��z�vb�ۭ�����؁��N�Tި4�ȂS �D��3&��6s�
��9$_߸Q��D���jߧ�����w����5�F�}T��`�M[X���}k`@ˀ+��6��xf�E��#�΅U&�o6['=�o7��?���F���o��_u�3 �A�&�箍A2C@"���>�ѭ�z�~�7��u��ug����ي)���8$L�Ǐ��N�ݙ}舧��귚�2���w �ABĄ&$A�����HQs��f{�f��h ��|wp���@`DH�h��nN�l��{���,C~����X^��+��m}�%ԃh�֕&l�C䉈s������-����ˋr��M�sjY�l����iIh����b�J��t����EM=ݨ"����Р� 4�M��Hg��w�@oӊ�E�}�����r�骡6���6aP��h@�c�Ͻw���sB9�+b�r�۾1he�X�����Q[����@Y�9N���::�9B��#�n�^���=u�4kՐ��8#p����˽��e�74h;��&)�C%E��I��䰼�xs�75�8LQ�j3��+xUO_|�q���+?��3&xU���og�X�@�T�(�Gv��= ҥ�{�w����ŧ�ҥk�5T� ���4Hi@�j�	� ���B[r��h�����Uuˮ���v�۶a�4����ye5��~�k~_ER�7f\�̢#�����l�x�z=� AF��	����.]^�P���7v��Õ���U;dy���E�L".Y�tO��f���� l<�����r�ݿN�X)��d(�Gw{B���;Z����1�/�W.�7��2nai�1f��f|�}F,̎¢cM�yV�L9��w��pؚ���}u��
�DU��0��дE�>35���gmw�tk��,�I0��,m$jM&��B�˫�=��.B�F6�rAp�c>����#�vc�3˃fn؟9�{���?'a� ��ۑ�eE�Fs�a�����'˹��v�g��P�d���=�@�������nm��c���e~U�<=�x��:r�D�r$˂��8o� ̛�C������d�_8��y9��QF �(L�n����,g���w<+���;1��㙏��)Ȥ"8$L�ǝ�q�����˕����{�z�(٥�}�m#������� �o¨w�ӻ���+ԩa���t�7o�#��fB6���9T���������7�b�VT�"��@��T���%S��Tl��pI��x&F��VgD⨫�ۗRr��;�ڈ�K:i�;�=[��-n�n�l1;l\	��u��������v�lg�ݯV�\q�q�By�ݫ��=b�K�8ێ؛9E�ufW�Zϋ�n��a����O\L���>F�Д�c�l��n�V�p }��m�(�k��4s��͓h�Gh��TKŵ����\���'�:v���f�H����ݝ<v�G99˺�w1d�pg�m�l��{�=��p{��������m	����Ơ,x����ק]��3��2n�������W[��u][�93jc�4I�H�dj4[eK��z��o'�Y�������Y���>91�֗Xoʠ�(�M�.�v���އoO�EӤ�ښ����
��K���2H�e���G�x�&�����z���t~߾�7��	e���l��P��;�|�2�1���U��C9���ʵ��@)"�d��S�}�����w�.-Z��
�H,�.Wz���oSn&YQ�`�$�T�En��M���tS	Ý���Ά�u�X�������r�ڂ��f/���Ѥ;8��Z��p�"=s���<wu�{�̨)�"������U𭉾baVd7�ɬ���}JP�x�f��:����P�8:�ؚ��f��#��[���1]���'$���VU,y��X�o�^�`H�cbAf�;^$ŉ�h�x�[H�`�Y"�˛�.�;�u5���v��{x=�"
4��[#S��|S���w���{����Ma�N� Y��Q`"�	&�F�w�����]��qc;�ww7§������^�0Dр$��H]��4~��]n�� �|Sչ�7sE ���l�H"!2@J
>���뜅��3x�ueky����p���;X�g*�m�6h���� �����߽����5b��p����Xl�:�T!���U�t�$���w��ػ�Qd��p����.�������jŹV�6k|9���~�R�L�MlU�}�#kmR�y��^�����i���2��I9��MH�},�^���mK�q���ރ�Zraf�R+,*��۷�e%S�3�,8*�$��P�+�U���]��(�����I:h���q�u39����T0��U	[(�&f�cGux�����'_n�e��C��}����l�,h�h�d`�2�ז�7�Y�����xp��_7����|���kz�7���A�4R�C���[����s�ޝ���2�C�\�y���n��8g��4x�Σ�&U7���=
�&�f����H�pa%��<�R&�=.ի��;xz^[5r�^\��{X�Nv0�������F���F�YS�5�#2��z��,�Ǉܽ�f�ɗ$Xp��F��sNj5<��V:���F3')����޶��Rh��w5�;�{�� �!^�v�t����ho�)�/}���]�mh��M8�>�v��&$*����1�d��P�C;B޾�n�r�?+�ξ���{��+�b�Aw{'��;d:�?6|;�۲WQ�r��q!����-���y�f ߞ�����<�����1�}�@L��b6�b�]�s{�ni��..5�7�{�d-w�,	�Uy��ս�����Wv��s��+�:,'��Vu�鱮��F�
ɲ.�~EeXB�~�%뽚����q�]����
�N����N�%�wFrYR�\�r�h>z���h��˝�!dڛ�fM�R�̪�XGN���ͫoL"zg{P	�Qi@����}x&�:���ؽj��z����{N�L���*(�N�g��n�j[���ya^GMm��b5����{���(�>���v�0��]�4c�1��]�=���d=��W	��D�O =+�����3�ܧ�1�gzd��9����m[f-Ȼ�1XL+%�	��Q����)�=�x��Q\5-��N��j��3��u/F�*�y=�^2���|a���1�#�K�6��w���
l�u0y�O�+x$��C�HC��A��!�[�1i6�ޘ��]V%�Y�2!�_7�1�6�Gȯ��L��Y�	��ރ���'ɵA���;b�9l�Ɓ9J2K$)X[	$�Lâr}�X� =D�"ˑ���3����o���7y�� ":�3�	����dӕ�0��3[i˗h�7��'kc8��zAcVm�f=�� {tgo��Ԗ<�z��;L��}k^�B��vf���`h���3}����X׭kL�`��G�b���N�,�vb8��^01o�u���9������w��ॽ�j^��,�7H,A��O�='E���G{��v��g�@�MS7�wo;{(4��4f�]1�A黺�=2��og,|� 紩�q*��m+�<TI*�Ț&Ψ�cZv���RO��nZp^L�����Qz��P��&�X�bau� ���� ��B�aL��l�D�`�����؈ð��o��˛��#�<پ܌o��=+�Ǩ�[�����P�NqY�~q��,h�aR#!�����h��ʊ�*� 	�hjљ����8����)(�08�1�S#w|*���ë�<������~*o3�_|��_I�ʐI�b.)Rӱ�N����8ӥ�:"��nԊX��|נ�4H1�Y���*���;3Z����ت4B.�{Z	�RѺ�P5�4؂ᆋ̬H�~�VN黵�s5�=n����%����Zd��0�:[����Un���g3�y{w5���~���qq���H�i6�[���啓r������Ɯ���T��O-�	l�E1F���g����V���%ʧ�j�]U#�N�o8!G�WY���P�X��l�ȑ����!��FV���yQs;���ν�j��gI���f�� ���75����ػ����� hQ ѱ���])#k���絾��Lg��e�dH# �{�Y��ܷ�9�p��~�r�,g�uww5�����9��8����6y5큃q����z�N�;�;e���nnv��x�a�ce�H�-(vk�{�38���c���x
{n忠�]E$8������� =����ۚ���o'>Y�@n��z � f1q�+?.�fLg�˹ڨ��Z"�wT�4��ܡ�-؆�������$~^9-��f?�j�����]�H��sA2L���@0]:[��*�w����v����<$hF�'V�_��O���L��e�E�k���D3}<F��#!��.u�9��Q�2�v�qk8#� Z��a���_��6سֺ\�Σ�{0\,�2�DkGc���kl���{�;�S�]�R���b��E%�γ:pnq�v�7cc��8�����������d)᝶�:�sR��*��X��(Ƌ�g\�q��7l����l냧fŝ�6�ݸ�&ݽt-I��d��1�&�-�wG�l�� ��\��>�Ì��Ks�ٕڌpv
zy�$�بv[:�U�Y��w�x=��F������wx=�������5���H;7>�
��wE�e��e.d��H����zn-�q�Uu�(i�	BD�h}�3�2t�o�:C#g��詧�:"��>g�HI��p�n*i��]�����j�pUV>ߤ߮�"��������P�ݡ��˕�8"�����8����2�m�Yi4�3��"�h��ñ<24��"r5�b�	e2��PA�vf��z<;8�H�>*o/2�Ǣ;x���PK*��)@i�`��Rb{q����z�H;8$]�^��s�q��!�hCnh�P���e�����x�fC�#4�0hA�4Z��Ӯ {c	R4�#ʲ�Wl!۩����ɖ�`��&��3�q432��WGlq��Ky����Ջ2ZH.��	}w5
�39������w�b��V��C�&,IńR
I0��&��1\���Օ�����B����}b	HEH�ЍU.��F�wb���{�y��Y��_��Kx�l8D�-�5��Uy����4p��l�*f�=^lZ����r"�!��f=����o����{�����:�Vd~���`���r8I):�1,��|\!rݓ�7�ݝ��J��9��N��$��$CB(!����L�W�K3���� �����fcN�]J2�eG

F�/1�{���s�gk2rz��̙"��gh
��V=��FBq4$+v^O�}�l|�Ԫv�{�b�"Ĭֲ�NF�t��X�+�&��`L�9ѕ�M�8hm�\�r�4�s������;ʡ"�	��1�\�8�e%4��Y���y�Ũ��k����hѕ@P� ���|�����k���{���"1�̂\fV��UP��>;�=T�,�U:�C��̷�O�$��~l��µsm��%L�����f9����f;x��4鿢=�8n����ڑ��+�՜1NG�8K�����b�&�ؓL��@�	�Im�0Y�:}2�fa7��}g�<*�6�N�n�z�_p8�i�L��C�vw݇kw�@_��g�rm̝��uOVת�=�̧]fzPR(0�-�,c�|���/DJ�ފ�W�z1f>��/�n�r�zP�$�.��
o�۳2q�+d��b�y��	`�tn|'�s���o�%:����owA����Y�����V�{0i=�};p��oR��u�fq�����M��V`�l�+{����-r�����5T�4 ގu�sd�`�m��� h�y��<��� =�C��_O�f6��v�B��#��`����#)*e��*;��8=�goZ�=aO<�������q��ث-̰�>�&&Z���n�"�G{Ц�k�7f��$.3d��̬���u�=m���2���S� L���t�<�M4	L�0�	�H��[SK2��G����U�{(p�t�ӱ:������P���ֽ���9���fw�ͽ&��P�8P�I��Wg�����ވ��]�ElqS+�R��j���Fe�O/�b��:cme�ݬ��W7�S�cv��}ӳ7�ۭެ�7�>S���G���T�L�k�JD�Ł�J{m��]�� �u��N��v.-ک�8�uA�mo��;?z�ܱك���=(�{=�NG^8�rq�HD�N�7��^��Nm�v��8�;[���9굻`NKm�=l�@���gv�c��ۗwk�8e!�����ϵ3q���p��6�u����S��x]�i#a��WN.=��\�tMX �r�-�[�#Ӝ&�)�����޻x�����L+gq��6�;���}��,pI����vV	�^;lRZ��q��77]6�;����a�i����L��G����wSlh-�5����/;�F�����$L�D)P �x�-|^ 	�8��~<���^�L�o��ґ�)2ьDP��7��SK���{ќ}F����\�q� �E�Z�̕����<���W�c���#A]�˽��;���a�L �6(�J;�UG�{�lq�Kwk�T��n�hR�;RT�Q�c5dA$l����9���kcw�#���+n˷Q��[9-�7CE�6̬AG�˺��]�3^�#��GG	����M�B��d6��mݽ[^��h�n2�����1��@���԰]l����m�������g�w��5�a��㓬9�֫�蕋rD��u�Dl��^�t*;D�-��}zND�Ӟ���YŁ�B,)���@�H�F�D}�;��L��}绛"���@	�{�|�$M�$4�*7$7g���5Xә8*�ݫ��wo���~O��!�P��G2ohk�}������*e���sw���W��w+7"� ʂ�h��LEݤV��g�{ڳb�}�$L��n�»U�>$��ZiD,R^�m
�53��W=��f�yë�;z�;�˪�͙�4\��	n�s�������s��gG� ���Nt�$ԅI�ƋLfOrp�����]ى.���*���0v4�,8m�2�T{��$���y^��`v���N*�F'2~e���,���!UnI��U�'gn�v�r�zGK�*B��gɈ��Ew=���0)@�-|��=�޾�B���'�
Œa0�,�F�����s��ѻ]�?r%���!!�L��A��� �~���+��
���</�HJ�B6P�3�6&_DDvuTo�ǩ�$��n}�׸��âܨ�_K��&JGa�k�ײ�l7]�@�t-�[�^(�Ns���n绾5꣼�H+#~��Uh͆���]�bA �^f�uv� ��H>߮�}啙�T���W���
T6Μ'�G�g�L��X�{�¢�����I+�%[p`��2>��gt����Qϗ	u:�}��j��fb��@^�ڟ�Qح�jKV�J<s;cP�7w=M�YSt�������sZ�&���ѽ/�95o��E�vd��Q;b�@�ܼ��ek�r�x��`���T�3n��	�"�H2�H%�x<����J�Ѕ�`l�3'~�v�UC{:��Q9��6nN�"3:~L�0RH$���wSs�ΦWi4�l.������<�.+%��EDi���j-�a4���p��ő�g�tz"�{#�&N�%6m��pEӢM���B��յK��5꣜�H�=�Cs�&�
a�ۀC*���ۍp�!_Ϗ[�s�S�qd6R	�$�h�ܝ�����.�Gȁsq�?w�͉Y�{�P)�r(�,)��]]�O�a�陪Ń��?D����j@�$�ɼ��9�5����}`�3{։i���ka��s��[^�[��B�0W���w�����o-5�+~�Ѵ�޾}C2yc0�k0N�x,b&^a(�5A��A�ډ\�n�M+�s��e���S�/��,j,b��M�{"�v���U�*��N��V~]�d䴣�ԍ����4�0K/I�j�J�s+P
i(Y�1�im�;:�`i70�cp.��g{ˈ��g�����Z$E��c�{E�l��sr ^)�;4wg���΃|�Z}��~�c:K��5��*�(���jwԵ���(�w�K,ܰ�\Q�ӽ�J+���H���̚���Wt�í����9w>�M��j޺ ��3�=�:��������w�D�'00e>���v>�� ���XۘI���k�{rF,7��ǖ�4����c�zwY��5wh��(y�}÷;�t���I������Lފ�ݻ榖dߤ���#�����2�\��$�,n��6�0���*T�=cl���a�Sd1GY�w�����G��mc�gikE|^�"�'Pm��R��;Y�4"�W�6T������]ɽ�C��ER�<�EE����M4�`ś�#�x�68���������B���0�V���$�g�7Y �b2�)�Kk�R&-�:�'2��^5��V`j��1����UH�;�b�o��ed8���lͽٮ��.�JT��t9
�x�0�{�-�\٤�N�Ȩ���;��F�sj�]ټ�"�%�^��������=��r��n;���b���Q�ڌ{��;l��]ŴD ��g��Zl�t�sۮ�q��d�E��=�,cnp�o"�w8>uź�P�l�K���]��Sû{VwVL�k���*��rN8y���[,���vN�]�n���u���׭�v���k�����h+ux\��l].c7i9��;b�玷vD�'vz�lK�v9�^��,M:ۭ��O�6����1<4l���k�y��v�ƆS7t�;^y��Oln8�s��p
eW��KU��xz�b:;inn�)z5�o�An�L*%�:��8kuÓ۹�EN���c�������콄'�]�-���+�)�F�T�pl���[�T��q�W oWc��� �K�;��5vnmC���hz$�z���htj���$�j)4��.�!n�i����c8��v��ۭ�=��A�nL��on��Ͱ���Xnd�v͊�f70Z����24�Ϧ�!���㖷f�;�V���g���{�W�7>3���]����m�����>�{砍�lT�����kY�#ݳth &p]��kη�q�:x'��rs��[�ݦ��7B�*ux�i.���wUN�vmw[�������I.)&A�ڛr�M�8��*���vُ�*��n0Y��E�ݷN��՞ݸ���c��6�mt\Gջs\X�t���I�.�j���V�i�-��i���О�on�7v��p`lx�$�޹0k�-�p���Y8^v����#ڀ��5O���w�[�A��>^v�u��em��;]l��u�U�,'���s���7�q���C��v���=g������,�삏N!S�V�\�wh۩�8C���c��w�l��]�����ۭ`݄Ǟ�����˲�B{���5n�#���қ���e�:q��۲�;n7Hk8+';Tw<s��s�ϴs�;F�8^6}n�&7h;q��{Wg���s��X��{b�'�D�݆��r�.�VN�^���r<nG\��]�0�n�ٶy-�ۈΦ]ob�a�q����GU`��c�][�B�a�-���7���F�QlB���W2�&�x-<޾=4�W~�Qְ�?B0h���[��2V�W�.�{�A��«5�yzV���4"��pCM��/���O�D����n��-~H�D���л�M����aɮ��|���R|�_l�������7I�}Ju�p��c`��u�Q�7��-*��oD8���̋��Y͗�j�î� �|��@*т1���E���;�~Of�sG��w�������cGҙ�C��y��h>ǀ��!9z��"���8�͇"~W��l�:�a=��/���m�[OΖ3���:�}��ގ��xcؕC5a��hдC�ͻu�\�XMLkw ��b'�o��F�؎�?AQ���{eSZ����+���R:����sڨx:3N��� ���#��),�-hk��d~P �� 2u'뵊	S6 �d,���5$W�MI@��@�/[���n�J�0�6��7���2_=��*A�m��bsF��Q�T�.48S@	.wW�[�$�_w����j����_s�!l�Q&4n�Z#�og�����������Yٴ7;F���RZ]�:-���0��x>Q�w&�5a�:b�!��ʡ�l �h�7h�P�=�8��8�E�h�p�ms�!Ro.�����JUn^�:tT+�yg� �׀�1��e=8<4�����\��y�pc>*<� +����7e���\uNWU�M�Kk�xNۋ�Y1��Gl�&��@fz��4v����
;��~����������n���(����s����}�Wi�귭ǭv�����㋮8;���j���Z�wc�p�lp�!�"��pcc-�s�������y�5��n�I������u>��n3�x�2T�7fu�L^��;��m���υ޼�^z�����/�rĐ� F��Q�д"�oj:�A�8�)ڎ˸�\�۶;�7K���P�y8��B�&FˌJ	$L��Ύ��;���9��
��.��'��{��R��$RF�f����?s�^�#����Y�>��-�
m��h�TJ�#�kN����'8%9�$��g�(�E��3�3�@�։��ٟ��5��G\wU}�o2ZM$���,Зz=9�(����o���́���쟼΢��ěv���	�9z�\���!ux��i�9�f(��-u��wU�̓��k�~u��$xBDf(�0�K�
%��}�#�U\�l���9aH��\ư61j��&�.�U�8�.+�dDU� ��� ɋ1�S����mڌ�/�1b:7�'�CL$��P�3�CgV�V�u]�-�tUd��]O��b)D��|�?S�N����jsQ��������m"H� �<� 7���\\�~йv�*�ӫ�5.��W_��5$(��{��Y�;���8�}n����]���<��h��a����19�y/N���r�L�8��㧧t�5���s��I�Ĕ��\:���o8���\#�@H�1���� (mL�	�*�ޗ~A��Wk��w��}����N �)�S��.�xBEݹ��
m��|��P(+��:99���'_v'�(g~���l������\��w����$��T߼����/?\����3��ƹ�dQp�H9�8��.{Q?=1y*I�iM�&�!6A!��gj�}|�Ǚ߂�c�>���Р���ȷ�6R	�2���
��}�����[���%N�=4�x��o�M���q�tӰ�7Y΁2nՠ��Nu�CQ��)@��a�P����^^�N�7_�k=�=s��3��&AAt��[�=�mؕ?a2��J�U7�v���J���3�_y�����&_DD͕$���?^QI�M��h�TR���;�>�w˺�tBYY��i(҈��)�NF;�\,�����7�����Rq��w�����֑�q�Ơ�fC<p���q����W����\�����y���u��L��Dc�d}�M�Q4�3����J�U1�>H�ާ�&Oȕ;�L������?��'�j��s�zNvA�7<�5�g��� ݙ莺�X��m��"#[K+V1�z����)~Kõ�n�Brݓ�<��(�A(5G�c�ު���e�˹S�N��G�Xpa��"\ �4k>'�|cvTϣD7s�d�lL�{�q>�0�IcY��@qOy�OHɦ^z=�?ES�Ȕ���0@Q�ĵ��瘽T:�я9�껙纩�/����Q~s��q���|b��wD'�V�ڒs([�n&��p���(�~	y���{m�٢�E�n`����-�ýu�%�cH"`��4Q0[�Y�ӵ�2=ol���˶�s[�O�K�(�=睡�v����N����냄��Əm'	����ѿϷ;����|�p��>d���'9�N�[v��.�q�"C]����F�y�\G.t�F&�宺׮�w'u��'T���=�[��۱��wl���nwi��$a� 8v뇫N8xS[�)5�f�{&�ѝooi��p�q.�s����x�7�;� �`:/��ߜ�M�b�k���/�cI�r�]c��H���q��#�RZ*'�E�@,��O2�șg��P���ï1~�2e�R"�n)V��3�z"o�r�D���Y�S����,5)��p�Pf_��Q+y��cދ��z%N��2��ti)��)�S��j�tp�m�H嬓;g��UOz9GI�i^��6�M�Bl�Cn�<sbT��s�ՙ7Ͻy1%�]�5@n���c~������q�	G+w2'���Pm��̯������=9zUí�u�h��m.�YB����|>��e���&U~F/ȏE����J����aj����:�
�87��eu���t,n��S�͌�ndF�%�4���F����:�r�Ţ�ټ9J64�^s:��l;ٝ�2�YOTu柚îr���ηJ�{��E�'��6���Wã�w�~��qXq��H���ߣ�W�z""rΙU�u)��� �l��b'�!D.���^CSj�<��W��F��)(e�[��3�t���{�P ��A�G���G���Co<<���S����{`��ջ&w [r�V�h*�r<]�y��(�z�C��������G����2���y��-"��4��:#��G.�gFt59x&wރ�=��)�@�Ԏ���:ZK�~���M`�0=����X�uj��Y�8�����c7C�7�F�����B��N]qۖL���.�9�n��;9t��r�7���c����ڍܻr����}���9�<DA��UrN�K���0�(�A�� ��Fd�Nv�{��}���B�8�0(�E�Q1�y��7g�)p�w��.��e� <A^��!`��x^zŚ+�݌[�>���i9b�n�9k1�3W[h��� �(X�qw�Qӛ���S.�N��p����@,�G�w��R�ç��p��2I��"��o!�\d��)�p��]j�U3��m�����}��r&�`�B@�	�\UO{��è���o ��fn�|����g�(O�Y<����v�:r��屐Ȝ5��
����c%��
�W&���z�gEqWN$IU'�q#e��9��#zL��\��vˤϢ@�d	HQ4��Khy�\�o��M��)�S���'D$z=��v��U6tl�'��y���qd��(%�3��u�V�!�B������y�ͻc,f�&�lݧL��M�M�Jl�Za+��z%NY33Ϝy=@V��Ck>�4�r�M IѮ���*��z�p�2M��ʨ�͎�z�wi]	6`4�,"Sϗ�*tI�=@H������k�2{���a�%��K���>��;�*r�ٗ���r�i{ݯb����F�"3�}�~�>�=ooJ�ifUGꏕ�`=g�;3O������ :,��(&�{B?u]�uS<a��me�������V
ob��]U+c���*���2�d��߿��;d:w)Z'cc���ܯ7]5�[!�F�9��v2�v����������g�����Ϗ u�\p\r;�\�@u�Cc����oӳO%W\��+�&��ܘ��1�G��`��f��Yn3W9^Р�:��®̼p�'��6��^Ÿ��C[�<�s�M�:�0o;��b�ɮt�A�
�n^��2��8�m�>z��]���ԝM���8y�u��y�9;�c���'���If�#@�G/�-��&0�v�\��=����nGa�5R�J�/N����Swh�S)(e�[���{�2�V��ė�P<��j���|!r	BX!"�ٌ�]�&�w��oC����nt@�YE0
a�����3�#���u�7����	�S(�i�W{���3w��k㺥�����oF��'�	m-I�͉��z,�l�+>ު��o�_��g̒�d�$�G1�`���r���6Fsz�&�!+�\靭v���贈����񯉬��+2""w�z'w>E4�f���Ϲΰ����o��6Yܽ��f�y���x#�;�sz[�&�M9���=b�]p��s=�U�๪:W`e`�U(�M����t�[-Qۊ���C/��VE�6�L��YU�8�����=�h'�_x��`���Ϗ3�y�U����@��T3��@i� �JMĿ�܏���=Ҁ���{ޭ�#>�bhL&D#Ґfir2z*����}��F��DD|r:02���0��s� �NY�3ϸ�;nnr摶к.[c�\����	,��[2�E0�t�����wF���r�F�*����i�I�Im�KI��R�خ�D]�t�����k�+�O�
e��z���~h�h��s��N�fʛ��v:�r`�}|f\����m�$z	�F��6���+ک��?4�}�t�}�M#{�ߺ9�Τl=�/���6AH�]N>��a眝"&FN-��ixDp����v���W�	��ˏ����)�:��Ш�HZ�f\bKv�qv�[3�v^��V����A�W�/�c��Xv*���*mZȬy�"�J���+�Nm��ȫx��\wU`��ra���|�edd��n�Y�Z�mi3G$�U�6�nl�nhꍵ1�goK���!�l8��5��r7��}⇐�p�32��[}t$w����1�ü����`���=-ma�ڌ�J�,�Y8��K�9"R6�;v'M.0Yg�zܯHЛ�7}�駵�Z�ݡ�A��ޞ-!97&p�w�^����M�{��*'k�2{ؗ����>>��w8NM������b�["�x�+N���-^ˎ�E�`{��A�U�2�5��|j�5����w3�co2����臆����C7(+��qŃw`���N䩧�]�xҕ��?{ΫrN�L�� 
p(���ؽ3P�[2�����k��bO����X16�˨�-�h���ޯ¼�Gw�����ʗ�{I�V������鶹��QWs�P˃%�m	U/1���R/��#��Nj��/FdPUA��ۢ�*���Ov���+4���xz+���l��8\��vA����u�ng N2�7E|7|�Bs�6��'�m�R(T��ϺEh�B7{�
���4��
�`�zR��޷�y����yL�X��� �6�6n��p�c!��H��}$��c/�*n5�9X��
`K�0/wk]Ogn���8	��鞐n�!��`�Í\�|�? � `R̓g��׺��?n�b��7*`~P�M�{{#.���}�n���]�+��.w�fA��y�;vѳ.%��w��]�|���S�/d�
�N;�3�ǽ���[K *�GI����u�+����j6Y�۔N6aapH1�sM;Q7�����@ʢ�r:}�l�.������.�����KQBÒn?�C,�Rz���0(�\°k SD_C���;v	����E�g<#̋i����{r�5oP:oy�a��n���5m�ٍr�{��KJ"��ͣ��1E�����ù�?8�^�N��]g4;Z��h��ל�#դ	�wk/9��;��4 4�]��\��'�w�vNq�a֭�d:�njاqf#�xj�B%һ|w�ow�����%$ɺ۸��X��1@��w3_���r���i�!�W�p��P%t��
9����.oQ��7G}�����}ݖoeP�)�[�i>I���RK.�thf -ђP��9�ѯ�0l�B��`��X��g!��xa�:��˭m�hZd�g[c���s���`/C�#�z[�բ�!��
h�6���S�� ��mU�����wO}��^<t`�Ӎ���nC�l�`�''f�۰*��q��:�J5f�jy���h�]�ډ	�c�=�8o�L�#7�:����"�iY�����ҹ2q��Ib�#���4����3;�V��C��&XS1����>�����B���3r���ݭ����bEӒ&�e������wo�+�pn���]��3�dĺ(�w�)mVn��b�팋��1m�t�f�763�6��0=���E�Ӻ�Q��J��y�]�����9�T��l���$o�L��x�����$��.o�{w� oY�r�t�/�wʪ#����D(�ە��1�*I��G�U��S9��'�{[)"	�Sf�]脖p-�n:����ꩩYOzY��}5**��T@���n2�T�ჸrSSRR�{�M�w����@�����`D�K�\��F���BݜS��--��\��РDFa �"�@3��;Ky��"�܁6efs���U}���W�{�Z8���%2�\$0ш2̂��un�{��z�q4�j8�A�lsR�dg��;L�%ݞ���F�fʒmf�
�sbfs���{�D�6�0���^�OP�mpu]�s疻��+3� �����.`28
��������E{>�qvp�s�1.r$�ߪ8m#fz���fb��H��C���rǚfc>���2�,%�Zn*�>�12~��k��ݒv8�9jd�~����Q��\�|MB��Nt�ҷ��v�M�)n��-ۦ��C�l�v��V�:������H��i]]y���P/�f1�t-�e�֘�oa@e0I��b��>����'�'���7]4>x�݇�:E���zx��.EI�u�����8�� �k�m�xm�7<v�%�.�]��	o�&�nFG�����d�۬��S����F�c'nw]t�m��i.K.�λ�� �I"�m��.Mգ-���E!���4���qNН7<�L�zC�4����G&�I�zu�K=gkGb.t���]w�Ww��}\Ƣ�]ݮ�?����ɮ����u�}jpq�mq�r;�ɬi�����W;���P����C����d"[����F���ʫFltz*�7���ϖ�(�e0�a8N�r7��
f�ɾ��z��-:#ԑ�B�p�#Q���H�:y�w7�Z7}���;����:PqaH�؆���-�ű�<�Y��ZW	
R�{���z#�W����w�@�a�L$�dfb���sI}�UNǙ������kw_@���"�OXs'����\��=Vf�5�|��G�F�3z�ڔkg�YvGh��������7:�����#� n�+ý�x߽O�M��I�KjWx�K��4+��(d�r���*��$���P�E�ny�{w6yz�l��7����L�M<4v�W������gT���>;�RD�gu���w�?^�ğm͍���)�@f��Ϲ�kw_������
Y�>��H26m�	^�k{�"���ݧ]�z�;Jf�#2�|2F��pBM�bI���=S�AJZ���֍~k��+͢:�|�A��H�0F
�4���S=�z��J��W�XV�
R�DB������k9���]��x�8�n�n�ׁ���[�(Q�ת�D���֧�]�گ�߿��L�{:*�|��?����J�C�`�Q��m(����kw�Wӊt�v��;��>��DT�����8L�,��d$.�|��S�H�l����Ѓ}'��s���2љ��,1�����Zv���8���P�r�3�
ap\��WT���We<�f��8P<�*r]�zndoތQ��f���q�]�}|z�y��߻�=��e}�К2�b@D����I��z}{�=���y|9��(OC޼�Ї{�Y�ah��ǚ�j%ڠ3����8V�/�7]��{��?|RM���+���׀�&h��J�[�j�璯]�#c,-n�l�RD�D�P���Fd�������ŧi�$r7���3)/��̣0��i'�]��Q���6s{����]Ǽ���������0�rD�����J���̭�y�}�=�kJ���#�O�rE���%F����.���"�������%�����ª���`JN����wn��I�x�ø�4Og0���'��rC��x)��bQ9'V���UW^\	�ԉ͎�0\H���P����`a��^n�G��i(�0���Y��=׵��ヴU$s��n��k���͌��
��ɸ���T��˵�d�׌��s�h��3�{M0A@��a�L��de�?���wI.ۻ��\�3$�{�kw_�=v�A��B�H�o_ޏEfFϛj�EEU??.d�P�{ӤyGqڊFZ�����U���wލ��M��#��sw�]��p£��H�̞�s�:7q���uI��3���T{�f8$�$�4!�����͕Ę�EgF��f�S62f�rqb����F""�����6��ubh��j1�&��;�C%�J��坋7I-����=w.��+v���v_z�x��P��-�j�""�C����÷s�l�lpjc��z�]��y�ˋ]:BLN�7�s�������c����<N�T�>�pb�K�8�x�k���v�S�nF��#h�	�8n�0�=��E۰<��[���xロ�q�ۊ9ٵE�5����dٜ(��u���ܯ�غՄ덑lwL�.d�n�i��u��@Ϩ|�*p�j4�7'W5z�r�FvZ��q��x�w^.��r6+��^/�w�����Wi1��Y�ȷ[c)؊Ͳ\e�Y��'br8:7jd�f�fE��i=����w������k�z#3�])J]�g����pR �w{��S�w7xtfc���L��×� L�G9�
�����n<�����n����G�DSx�7��5y#��E���I���ʻ��y����sI��3O1����x�n�+�к�1 !��FbX��Ýٻ�<������e}�̗���?�������Z;W!Lɋ�Krq��P��1r��7nz�Z���K���ɴ��T$2C��,Y������4W��b���
���ol����J(c��w�3��ob�Wi�_Ӳ��Y)�����Y}q:fQԀ���sf�o8N��n9��2e��@V�5���+�)lm$6�Q�W�fw�]Y�/rgX�����z�.�˗�[���㷷���w��΁Cd�矢h�32�p��v�|�)Z�ͷ��f}��Y�QUK��2�*i�L'	�B�������Ԧm��T�f��UtDC��h�H���2�>�H�Ql��.���
��v�߇S�H�l���C��ZD4K�t�m�,�'k�v5���s�ص=kVtq��h#yi�2�-60��Zj�.��X�9&R��f���d�}��J��I!���PF[F�esǹ<Vl�����s��%٢�U��y��(#�H"A�d�Z�����l�fcU��=��:�����2�Q�V�;��ԥB��A�����Δ�����ܩ�g�7�uC"յ�a�s`yS\Mհs�+^Xxft��>:��w]77;�77K2���&1�&F1C�=�_u���K������Hi"-{� O�J�K��z��-I��y�F�;���E(L&Se��H?UR��QUK�z �����;%L���Wj��G�q1����!���=��bl�L�&��K��i�/[u�k��E�Vh�R�ŭ1c}��߻��}���3+�y�ݿ��ވ����TEӦ����՚P	$HF8A�ٟP㳫3�gz�Vd��,LY�4�Ww�9t����ov{�Y���#�:*���q�Z
84�1��Ap��)"Jj�lzk�R�f�)������E��Gh������d�L���]���CӤ��,'v��~��ʠ�돧��]�3���̘��ao-Y����싺.�/�\FL��wk�
����y�nhF\�o;�]#�N������;>�H�q@�F4q�/�<�~��ݼ�}o>|�ջ|M
��g��WA��Ji�]O;q	���'Z4e1*�\���d�=�b뺢A�q�ڷ�?t�m���fd��� 7ol�x�f��;:C�(�`d�#dkݟ_{o|(|�~�/�N��f�*m��]�DVd����*�Cl�uo�TES�h�w]��]�����9ou����!�dC��7��kN��?�ٷ�>����'q�n�l/��T�L�&Aۺ����\�{�w�kuk�>�R�4)ӯ�����o���$��		!$������3����r�ڶ��ջU[k�m��F�j�ڨ�����U����V�Q�X�6��kTkE��m����ײ�ګ�V�V�X�m���E�m�Ƶh�Z-mE�ѫmcmm�6ն�Ŷ��,$������������r'�BI �E�-��_���_����!���y��~��h�����~��a����V�~_�?i��?�$��_��0�������@$�l$��D�P~!�������~���	$���g�?���ܣ��y���������ʷ�m�T�SYU5���k*�Y��ͪԥl�T�m-5����miU�ZU��5��ҭ�Z[lڥj�Zj�kJ�V�m�kJ�mim����֛jmim�֕Y��ښ��ҪUe�6��Ҭ��m�ZV�֛m6��Ҷ��mi���-���ڛZZ�֛Zmi��kJ�VͶͭ-����ͭ6�mi�ͭ-��R�6�j��V�kMk6��f֛m���SkMm�֖՛Zj�j�թ�����MmSV�kJ�kT��m����imJ�Mlڬ�KU�Tճ[-������-���R�S[J[R��R�6ͭ���-i�em+T�ҵM�-�[R�J�����զ֛V�ZV�miZ�ڛU�Եl��m�mimY���f֕�6��Ҷ���Zkm6�����kM�6�-i�����SkJ�6�մ�Ҷ�kK[M�6�f֕m�Zm��T�ڕiV���kl�ҵjmi��MjV�MjkmSkJ�i��m�mi��6���fֳ֖V����kkJ٭��5��Z[jmikR֛m�jmjV��Ke�M�5�m�kf֖�6�֩��V�����ҵ�mKV�֛Z�kMkl�Sj�5�kjj���5����T��ͭ5V�ZU���ڥ�-T��kf֕Sm�ikM��Ҫmim�i�*ҩ��٪��MSkM�ٶU��M�-�5�6R�5)YJ��Si�JjST�ҕ+e�kMM�6V��kKf֚�֚�����ZZ�kMk6����եm6�kMl��SkJ�֕-iT��i��M�)��J�ٵ��Zl�ҕie�4���ZSkF�)��f֓kI����Zɵ���MT��M�%m)��6��kK6���mi6��Zf֍�&֋[2����6��ZMZJ�S)���M�3VM�)mi�֙kL�ɵ����֓jSZ�V���M�%��R�S6�m�����6�mi5i�ѵ)VR�J1JR���M�֓j�Z����E��m��RU�mhգj�Z+h��j�f����mh��Z�6�V�mh��UQmi�W[mͭ��V�kF֍�Z-h�RmZ�[Rm��kj�ƶ���3mFڵ&ڛ-S*��S6ԛjfڔ�*V�6ԛjM�)���Ԧ�&�)��mMJ��mMR�ZP�?3���~��� ��H� ���]?�d����p�O���������ܯ韉����$��O�~�������0�L~@	$���"j�	$��� @$��4�~�_��`ih�Pz��F �@
�G��������@ I?^��c�w���t~_�8���K0 �I�{�� I?����JS�?�8��1��xg����|J��:��� �Iz]�bi?�g�:s]9�� @$�~��^3��� �I$��/��������?���Ɋ
�2��ʡuP�n�������?��~��2�=�          +w�   �    ��� ��(R� 
 Q�� ��p����N��l<wr����Gln.ue��"(w���]��{T��.���^��it�-�ݳ�O| �q�|������U�<;U:kQZ�����(Tݱl/���V�*�v�aG�<t �8w�t>�l(}�T^ϻ����v��J)v5��w|zM�UU���i�����|��  `ؼ����A�w��c�Zroνi�T.�z��M׮��̏�[j֮��UoA@ �{α�f6��3v�5���d
�u���{u�fow,v�}��ֵ�     ��*�       �~L$�T��     ��UISɪ�0�d� ��0�& j{E*�� �     i�5�� �     D����	�(�zi�Ѡ�	�z�S��>eWEP(~��*��������DU�#����?���I �����/�iO��� ��@�@� U@�w�~S��'�ʀ����}��?6�����?S1�?�X�>�E�q����YԚ��dsw_�x������-��;� �z�ǫhe��Z���=��8 �
��ؗ=F���uS��F�o���H�x��<�!n��"՝�S���:�{��w���ouX�	1�wF�[�XpǓ��;g4�x�� ��1�\���@�!�UBp��� �����m�ptD|��nW���ݝ��8aH1պ�Z`$7{"}�vk�5ւ��������Ր�\���t�se�//<�P9n�۰��9˓���x�l��TXs_2��56�w�m|�p��\n�zH��2�� ^�sw7Q@w�s�^��Ň������5+l޸��b �	��Uŧ����N��Q���_6۸u���MC#�wdۢ�u5G[�UM�H�M|O"4�cI	3�\���Lܗx���Ky���K��&�;�%ݒ���5��dD+�Y�L�WV��N��5�i#s�[�����ڪ$�-\X]�zc�3��@/��Eñ
�u�j�r�!΅�	���2����ڔ�n�p8��8]كz�������d�,(���Ov���/]���1�J�7L�wl�\�q;3{p5����:W΍፶VI��7�y$'y,�< �{�"��;r>0�h�8�iՒ�v��{ۏ`��d�]z1�dz2�����@Ʌ^o�؜ �u\3�{ůgJ����;2vl�Q���oEQ�΅�9���+jƦ��"m	 ¬�_0αŋ*�9�w�!� �~W���B�PN�[� :y!��uoUt�=�fǛnڹն\�c�Z��SI-&
��#��1-�Ԧ����;N�u��̰=��b���&o���}ǗW�9��v7r!V�bf���J����*����B/
�mdK� {��E80��d���2�%�L�����]�1�n���7��ߟW7����添n�����Jg�n\�n��5�^�AZ����:�J3r]SR��X�m�$b��7LO�:"e�N��v`��j䝺��킵��C��Ů��$�J3�;�r%�ŧsx�`���6��;F�[�+k�BYϜWb�`�t<8���&7�LD,�n�۷��΃�6@r^s[�ָ{�#Y�h���Y5pc�tPz�&wr�T����%�;&I~G}ۆf��}ҙ�-تc�tOP�)x�P��[:A�M]͹# �wm۽�
�2ݷ��[�����m6�x���,����4gq}nɔ;�r�iw{���	�t�(�F�]�#v7��'yѕ�0Ë��٫R)M:�����b��V�ې�U��q�i�Իp����myՃ������.�1�\3A�&\	�\y+u��8fY�wm�լf�S���ۜk��-�^���gc�ka�p�{,�HÓ�w�y�sC&Hܽ�\M]��`]-�i���n�y4. �0: ���+��/sZ6��>@vv-����L/.l���u��:� IMܧ_�P����|5e��k��s��se:��ugK�	����.C�z�j���i�y
4YYG	�dZX<�3��lD\C�"�nee���4��1�lkx7@���Ƶ̴W>����B�uS*K}Ŗ�@��{�<=mZ�q�dػV�7�`Su�,�g,��ˤ���B�'^��l�׈d��q�=��"㊩�ݦ����?8�:^�x����!�:9a؄�&�79E)��U�0�"����#R%��P8�i<=Ě�t�� V"��,Y�zE8.�18�z�B䨀���(�n��U������p⠫%�.n.�7C��Õv]�>j��K�.�.�K�S��RG���3�>]^���;7�\�U�n-:8<.L|�^���yv��<{�Jq3�> E��p��镁��a9(�nwN޸w��l�
؄I��H�h�p�89EA�`rg]퉽�ǺY�:N*����8@�&E��DZ˒�԰�"��2��VP�=Z�ȂOvQ�} �ol'Ӡ��w��[oOt�Y&�&֐o5s'{c����~���G����~��v4h��c�����*b�����'�Y�*(:�������Y��(0�V�=��:ۈ�����M�:�����5����uU��Q�i�;&T��C(����8��-�z��%N7�[q{%+��؞��\v.x9�3�K��5μ*�G�o��u��:�Ԯhv��۳��ur�qp�K
oc����1�p�[���.8�v;���a�ke��tt�mwn��rv��5�N�f�͌�,ێ[��;-��מ�:�Gg��ۯn��U�����3tv4.�[=�v�.�p���c�������ώ�^��tk�-`3u�gĚNj;�Y��Hq<�os�c|�u����Z�GM���8�ѳ��{X�w�n����-s�8�o%Kv6�h:��;s�/q�����͵�r�5�۰��<ԣA	ݍu����i{�ՠ;l��7��n�|�!xw�4���n�omk���=�M�7�wm%�׉ې�%�����1vﾯ�~[����^�p[��A���tvs�蠛[�=e�;<�jt�s�:��y�u6�N(�';���g��;����n�\-t���8�ŷ��=f�E�4�M�q�<&��G's��g�clu��S,nJ���A�i��z�ɵ�r�3=�k;@v.��A�����ۣ��/O7�\��ϝ��t��o ��۶�Mn(9��Q�=ʨ��vG<�{Cs�C�cU�:��8{Hmg�Qɵ�k��m��.�;���:�S]nW�js���f���0�&N��A���;@l���]1�k�7E�J|s�yy�
���Nwm=(�>3 )C�g��N�������l�3k�7h��_�u�3��݉q{G=��I�υ4�ب����`�b-)��ʷ�Dq�Y��M�l��lOl�˞�M9K=z�W�=���P�����:�'��rǝc'[X��lp�m�v���N{�4�w gmӍ��V�MحΝ�����v�;]u��{A�{v79�{����s������	r�;S*q�R�m�;�Ӵ\��@��ػ<��쎭�������Lm�e5�9Uc���]��^`�٣�wn�n�9�Qԗ��i��e���Cѭ���1�񻢶�5�pj�� �q�t=��d�c�<<�y�O��`���7��Ƨ1(���5<�=�<Bm�*n��&�z�8�Q���V6���ܦ�ݣ�ۚ�Ֆq���V�\C��:�&�!۝�X=�˼�Z:�=lS��{Y�$�n��1����c׆��KͰ���#jz�ɵ�����8;s`����Ҷ�0q�eV�=�C�9�,�-)Ը�xU���)��c+9��+)!`�L
�����?4k7=�v`PN2���?;v��F��h��V�-��,j�lf����kE�*\+�Zú,=���Ul����_2�ׂbk��Z��ssqWSq����m��*v��u0�ik�u�!�����M�S�B�s& r0$����rȖ㳈�h�./���~|���㫳�1�ݜh��ȅ����@�}��Z��!��, >ѫ���b��/�����I~C�u��W�4�2+l;�UZ�H[X7,Jx7��ו��)�O�ga�C��0�q�G������}(�V�D+�7�[�ܹ��{LF��^�`�sj��<>�tA~y�H���N�-�z�.�u���=�y��Qq���0 �޼��.��Whf����g�>���I�[��3}k!��	ȇ�w'i�����[#]±���Ӻ�z,����o�ְz�#��_H����
���o�3���nN�nA�5j��Q�{\ː�M.E����o�H�JD��O�7�u�cm�9�:z�������nR����U��Ń%'s��|��սg�����'Ծ�����/o��.=�W5�	�����X����;u��C�43X7��b��=����Fo��|�{騾���G]��/M�ё-�	�|	ٹ�6�+��z�-ry��i�^}vy_n\�zD�e4Ǳ�FF�Z<!LgfɾZ�]���̙j�ꃬ���v�}�&y�O����	ʎXk�U��z��Q��R�.�W�4g=��=א8�
;rLE��.9�
��f�n��@yd���R�|�������:S.ʭ�9�f=�� k��Ӥ�닻
P28���ǥg��/@��j��g*�WҞp���=��t�Yl���}���QH�4'�7��������[�7$Bj�wx��ڸ}٪� ��6p�7Rx�3�e�H���p1��\�|�)�mv���k7�2uD_��efW�U��x&w�r��ͮ���Wq~#Wx�o����OQ�������#H��dE3[js��ěȽ[�6�ǐ�Ò��հ����ĭf�6�CV�u�=�#���@3��A�a�D<����ui7�='����Z���gk�k���d>���^Oo��<�P�z}�݌2�=��}�����<8�����|�}��ߛ巶x4�t�	T�Ek��Խ{�'�ѷA�dZ��5[��%E	���s� x�'�ᇥ�{ٸ�@ݠ�շ�Nݦ��U0�i�o$��Zk{�������h�ge�2�����v����Ye����ڹ��^�3n���o ا��hcT;��_�_: �.w�y��`�m����C̬��{�ϱ��q����v�ڪoD0Anr6Wu���r��q;T#Ӻ��{���L����鋣\�v����zcn��86Q!�u3q�:�~a�%����^�-ݝ�W���![��j����#=�8Y�U��m�21�dFcT�9g%�S��ùD�xby�yv�E�1���ϼt�D����޶������Ծ==�]����׻�ٻb��3���#2ዺ"�]��H���� ��8���^^����O8�8���y��f���]^�{N�p�9�9�:(��ݾ<�]#�wgc����9wu�k��,�Ef1x��f2��2��u�0�M[ա�2|.��WT��}�9��V���.�ӻ�gx��{�W�#K�ǟ\EO�׳S�k�gEC}��19� �����3�m��<�ռ�|[��N�ƺ��~�{��q tՁx����2o_n,cZ��K���w�f)�ɞ���[�ёi��,RD�� �I���t��\���}�i�<�;�~v��%�`����G��E`�Z`�^ο���A�D��>ާ��@(�Y^:'����9g73G4F��g���nI����]0��E�K�!���u�;V!��t��,u�;�H����[=���K�v���{��~�nd��&�dX��"�g��x��/�^�2F�cnJ�]��=�Ǩ�|�w�Ս0��|�1i��+�]�W��gw<O
�ZLC٩��T�F�w� #@��<t`�Y�{�91�{�eBa���r+7P��Cւ����=���8y��?*��ǻ�ݽˢeTz��	�[���}�=�F�Z�g���N�:nz�-�v{��ږ0j9q�6i���4�
�v˨�Q�3�N�V��6b���שE��˲oe��N�3=�L��O �
��H��~jo�Q}p�L�X������2~�>
�%Bm��蜹�+����m��S�o8���ϣn6�k��(�)��s��n7�;�����ueW�Ǌ�9km�q�=���8�{w+6^#�Oc=�<����-�����:��'`�۠��]�l2nn8qs��m�ir�7����=��`�ç9���[axx<�՞Ŷ����\n��Y�U���קr��y8��nWj����h뜺��y�t��kt����n�iݻq�z�gkv�޽�pO:�v�Dۮ<[������x���SG�7=cG0ۛQ��[�Susv�0���$�ִ�*��������j�;Mak�y����-.�����w�NN��dz]Z*#ZR�w_M˄�Ah�;vb�f�H�;��,�{�[M2.�i�jD��qI���N,�Ps���=������}9�o������qw��=��E03_�Ǟ&ת�MC���)��)�10�1qDBڍlf���/�m��9qX�-��>ϳ��I�J�d��N]�
	%	�qU�#1���d=��ݐ��ܞŹ����Yz���5��Ѻ�]e����݌��u�f�c����H�;l��<�e��=�vf"ȴ���|��w�@�a��2HF�&UɃ5�B8 �"~�'ז�}=�]��� ���,�`�r�!�<��̧�A7�'LI+WD$���^�mT��w��[���n,��TF�R�Z}���q��i��3]'8D�t'���O��k|��Q��B� �	� *��

B�h��i�5�j�X�����0�{��?2&"�����P^�v=7��qU��"��,r�9�M�}�=�+�V7֦��0�)��E��KJ��c������k�˜f�(�gE�pN!�t��r��A��A�!	�H�TB<xY�]Z;N3�~䟅c|���r�}k�^þ�$�Q8�Y*X9-H�����ϫ�`�Sy�/=�Ȧޣ�T�`."�29t���ku1HmL��4ۚ�88��؋GWE��(�J�S��Hm����} �|��E�^"<��Mm;m	]�R�W���DA;�����Cy�3���(�zO�aI�VEV�n��j�i�^(�ϔ�-9�R��K2���34N�q�s�j�լ�|7�9�Y�z�%�b(|�=Z�]s湃���C;vz|��$=q�Ę!&���vq<n���v��b�j��D�ULhJ��&YڽFR�Y08�J���{��xu��b�ZP0uE �=��0h{a���nH�k�,�U�Cg�a��C5�<;/�s5��X�-,-���ʬZ類�5��?)�쏻���������-)^��ߘ��Ե��3� � �N� 44��$�M:c[��'��&�8I2�0���D89K��-&��]�@���dW���6ʁr�[����Đa�@}~GGݬ�!�����V��d�(�<؍�Ep�:�v�7+LF�L��"ey�q �4� �66�`x�JJ��o��E�]���Y�{�hᕽ�t̶:�n�!l����i��0�P������N�4d�T�3�j}�+ݑ��&ڃ�"��<�L����J��'WUe��j`��f���/��!��"�$�ŧ��T]>�6��k�ڙU�!Hf!$Ƀ���XI�a��F�	�n�j@6�t�9��<C�E�IX���x�ވS�o��ƈ�+Oj�p�sU;��E�w~�o�;��d���FS���k;umĂ�=�ݦm�6�u�lv�{t0gsϷnok����:�\.��Sl��6�C6�bBi��!��I�!
�&`�R�*Z����-5���շ�xF{J�R�t�^YK7��{+S \>�ڎ�$V�x�+Z^	UtmD:�+�YG�,�/d�a��o(O8�Ji4\U��-�2����I|'~����h��(@�I� @� 
5�_����\����E�Y�6cb�yO�m�N8������ae$"*�,+-�Ga����}'�Uڝ���5Q[_�=� �x^�X�e�ek�sq�-���pcGGkXj����;�5ݔJ�2��
��6snU���N��Dqר����G��bHY�މ9X̎
���S�Y7q�uz���=�·�Vqő����L��Z���g^��a��� �ɽ��ys��!��v����{l�=-��F�+li�u��G���۞*?�P����N�7@��{����8�5q�"6�\����K[�+���DVH�9�"
���� �����L��i�e�%��fO�	6Ad`C���nvo�0��U�Z�w�<��(��n�Y7gE��'��(=��qlI|5�x͔�&wz�H���5{N^L
̓s0�5�*�v�2���]奚n̴^ 7�)�Usܦ��q�<ݐ���&�-��0ȕ&j�Dۺ��WZ9VjA�Ჵ�O��ſ(���.b����Ήb<t\}��r�� �R�$e`1��BT/�g7[Ϊ�+��W�o�"����8'�@h��҅�c�8y T	�d ��%m�,r�-7�OsG�q�����BQ�ص�א��B��j�d^!��R��S� M����o������j591��$����C�Qd Lbi�Hm�I��lE���b���f2��g��J� 1���8��)*��	Y�,bʐ�k����ѽ��w������a\���k~�����b�a�^�~޽��8;{���X��|��z�<���G,#�����}�����5���s���x�X�I��B�	xn��r��ݩ���wXl�c�}�3�ȼ:�6j�WE�^��[�vY�\;b'�/���o`*`�&��%ƋDpnF��ʪ��)���Iƻ �zg�����3��r���mP�+3y��7�j��7�<�᪇�g���xW�d�s׋�}���J���|{S�@�!q۹agj�-=Ew���kܥ�J���z�tˈ*k���T��қ;���JS_P��7���o7��ii4!�m �	$:(f56�Wõ�BVg�9$����8,��d\UĒYj��U����G�@����\�<�#u=ͫ����n�(.�T��5�u�d�iLg�ޫ����0��s�ˬ�A+{�6�}��8�q�)��9n�i�4���碓o�|���HB^n��*�*��	�܈h3�����8���}9�&��WRU9����^B≸�W��V�%�<��铉.a,^5�v��w�*����G`�+����Ls����!X��'��O+9��D��h�g�^O�= �ٜ��="�]�L��E��m��xWT�BPS)�y$��]:vC�Z�����4'�+㌧�m�C,�G
�mu%�L����&v|���c����]�;<w���MD����'o��³��	�Ò���q	{����W�۵,�uS��I�v!h.�ܡ�����^}n>���a��S���2�(��:T��'-��(Z�
Q����L���B��1�.�vz���żoX�:�1�4���Z��{�����rM��Q,��4���\B��i�UR��Z�;�F,UU)�Y���q�z�*sw�����qPα�˷SK�D��=��,X���8�P�	��\b!C��9�$�����Mk�}��حM�[n�/ЊVo����{��YｭTp>߾=Y� [���Q�q�83o��0nHO"	'T��{���m�<�����Qf��7�/�]��L���):�����Tu'��
`�ɿ�K�n'$�siRC����*�*�=�[_"�V`|���"��=���UD��"�����l�����T��L*�s�L�ݯ���,z}��I]��۔�*Wb��z1�s�IoY��6��~���+J�IH�����-����l8�U)%/�3O��iu�uRR�6%)Rwx���y+�\XX���]��9)�c��W�	��#U�S�N��w쎨׶+*����4���И$����>|k]椸�����BK)�>�ҏ��6�t�UH��Jȫ�XŹ��p�̵��IjM���l���v�J��� �p�^������? �K����GB�-}�+��tn�'��ˑ[�N�����Oj��*�rC^�4���W����{j�%�|X�Ȼ��5�k<�Y��j�&���
8�C�s��&��*U�]��Z�HK�=�Ӆ��K�Ѿ;�eas���hbg��Y�LY�]W����l��U���u��d�1�A�W�(�f-�GW�هԏ-�Ð�^`0��ݢ�����=����;�w��̿Lg��n�y����D��uQ����#z.�т.uGn�˼Х�n����`�/b�,n`=�Q�z+kz� T�C������@̣M�U]��ZX�a�������[��ҧ���m[��ݷ���qʙ�&��[5�u�f�!��	��2�&9pg�9ڮY7Br���M�P6���..�7m�Z�0�T&L�l��n�����M.;g��Ʊ��ܽu[��ol98p�͊�w�ϥ�NT�=[pv�r]�Fy|��s�p�u�Ji1�������T�����'���ٹ�nm��Xݹ�S�=.���x�:�5^�u��ۂ������i���봡㝵e�-����EL�Df�AS��KeD-u�Ӱ�t��o��#߆��hɄ]_�Hb�3���^B�?[a�4���Q��������z|��O�Q�rx{��u7rmEV���yߖh��Io�ޡøD}���)8�<�{A=������|�[o=���{޲v�]G{o�c�e�f��cd,bq�e;L:�p"{���]ьA~c'�����@ɾq85P`T�i����_���o���<4]��.�wO�p햨�jڥQ�"�(�cr���׬ #�jFw'�m��c���l��E��\��TK�M.�iF��pw���"�����Gn۸�I�UH��.5޶?[�H�{�ޙ��M�{�x
��L�c�c2A^��]t�g}�4Uy�E=�7���+y�g��C��6��c� �������*W���72�{$o��*���,.�:����٭A�kWk;K�UI��n��;�{32>��BF�����a�W[ʚ4��z�mrq{�ח[Tʠ�

 D�����Vyw;GD�/&���pC>JR�0x9�Y ���ʗc� �����-�ߐ��]��e���� 0�,�X��O��h
��!KT�;�+3�,�͊K����[7�C-/G�|4z&埐G&���L�.i
�l�<Q����	A���їQ^�¡��EXe���B�,��9�O*��+�]g=������_��l�]-�$�=�yϾ��C�W��}�,��RH[��'�5p�,om��Ժ�j�if�)sS�=@���m�V�z>�Ӑ��͚|;e�Jf���4�8�	�K��g�k��_.����nc`�T-���m�c󌸸s�\����	A@R웳Y�i�'��� ʍ?b�O<$/�t5��nQe��T��mW2�=��d~9��"�zk3 ��R�TW��E����Z�oL�@/F4��*�K�֎��-�\T�7KZs޷�*�����h�~��$�ka��~ʻّ]Ӛ�J�QTB��X\�ʗ��M۵I�xzv�E"��Hcr�&쩲�7Z��6�s۴яv�S��	20�;g������ǃ�� a��nVd��E�A��U��L̶����� �Kf���b׃�	��'��X�f����3f������͔\,�8���}�Ȏ���~A oV�����Gڐn�����9}�[S�6o���f(zV��}p���*�]7�O-������z���:��Mm)��((D*�
�$�&&g~�7-������8��ޫa��������9������J���ڙ7F�a+�o��K>y#�6��ϫڵJ�,TN@2%8��������MLd6>��9f����zܳ��%53 F4�G���6onin|�F�"��{�����K�T�*�B@

�B����a��/\��7'���U�&kv����v���Yo����o�R�E8N}!ə
�䌠�ѣ�25.������%��X��C���LT���iH�3��ϡ�cI��L�D�e��;���%}waI��L�^g^��A�$b	!g�_o[��ˏ��K��r��i�g�B�%E��#����ƙ��Z�I��x��z��E7I}͝BǬ|�b�>J�2y����1G5W՞֎4̗/�~�f��.J7��[�,|�?O�C�ؾ(�j������k�R>����.����v���u�;Z��7����zz�Ǎ����6���`,k,��t��
;�%¾t� HPt (��PV���\VJ"��#��-���j�{�/��cg��r���}���#�h*E�]˖9��ɻ�b��}n��dNxc�7M���`�3���A%��wxZ�~+[N�ݕ�q)"+�3��.�RB�����|{T�/���};MENWMa7��oKp|��
���<d�!�0� FH����7��uf���#k�M���0��'�N� ����bf��)�Kk茇[,��2�����h�;���Җ��J�VQw�
W�����Z�/��?-��*��z����g��?%%�v��Ì�p���#Y�L�
�����a���B���='��N��3���2b�l�5`��M���7�羶����>�-``Z7ϼ���y ��;����d�;��_kY8(lS��6�z�2n�L�e�6L���n8��Ju*6q��6�Q�Sv�<%��ҳ7��.�]�����C�A�>:��v�^�[E����׻iH��WСMk��؍��26S���@+2F\Lۘ콌�
:��+�����gU�|dG\�1w����B��S�щ17Au���\P�8��u-�(�N�ږg6�e�@���A�1��e�;����+'�L|_�a���y}7|;�}���"r>#_)�����N"-#�`����Is���w���h�s�u�:GP1�Nܧ�B�ށ��S������I�5f�t�D��^^���P!�{6��okܟ8�5��?GƋ��z�����bx��b!}m�JD����!:)c����3-y�[�Ϯͷ�U�I���s]v�g;J������/ި�k\���n��	���C��T��3�L����L����;��0g<����7q8:\R<�� I>�� �%��k��{�M�2�j��ic}l�U_|�!�@�U�6��o�N\��%Y�*���@��A�O}���f.S�P��k�(}�x��͚C@�$9,��4`�K3m��s�'3�-� �O@�9^�zg+�Y��Ќ�٣��ݮޥ�v�ΥqJJ�U2P�*X۬-S`X�՞�J��b�����l���sκK�+�-�mb�u�����ppacM �h��Kc���	lDe���$��%��^X�f��}��c��=�`��fŽW�r��ХW�36�BGе#��)���?�ZO�@
���}�5�S�_z�k�R>����ȋ*���
�M�N��)s�6i_���ek>���_:��8P���$Ψ`뺽F�S��Rs�9ش�ӝ��2�$
��Sx���������Ĝ��Io�}g[59��A�U�qo�|��>�ۦ>���'�%����/e^�bq8ڱ��lDo�W9������"����r�<�^���o͇M�ܽ}a�Ssk�,Ϩw�C���|��z�OG��Є�PR �սٶ�]�{OW�W\���g��>�P�
���켙�&��>�v=I,��r�Y�xr�$y���ʼ>�f�h�n>[�*?r(
����Qp���Sv_&�������bU��'e�������v��ٜ芤-V��x
��y���ԉ�<�w+�3��R�ȝR����ɚɋ%("�z,K���3�>Qe��������1s�/��Q1v�G(�b�x�0�{�/�߃�g��߈��57���	ʍuP&�׼��`�]bE^�[T�Y�LltP��7i��X���\e^]��u q���\���7���9�n.|&�#�JIT�2*��i���������8�L��'Xs\����9�g����P\̀M��d^�E��=(��d7��[��N����/�ZE����ƩMrYn{k9^$��z�Щi�Ur�GB�!�AV,����{�'�9�Am��G�jt��H�F3�sl�E�g�'����8ٙ.F�u�j5'-�2|��ˇ�ke}�f)��T=���`F�`�����}U0��jࣈ�-��q̙2��ޱ�A}:��c���q ���F��,�M��\G��#L�6MrnQS���*�q�W�4��aT�yQu;��4�>�v��Me1����{�Ω|Ձ�'/��'�o��)�>���ٿ��m�����vo�6~C@N�
��ʕ�\ U0��Z��P���A����jf�Zč�+��\߾X��0�Ҁx|�bc#{��yS�\	��s3 ��PY?d\Ѷ���;-�J���4��c��Fʛ�U+��n�cعf��m����Pz��B��'�Ͻ��Sm�?cb��>l�k�8�G�D����J>��H�>0�6P��˳QtDcH�����<�8�O�Com��ʲ�o6 �^�Nwp�C٭yn���%��Y�<�fC�~��dȜ�Wsu�d\NN	OtN�ۃ]J7T�L��ٚ�"�ݞ�&�����q�"9Ti��ݦ*�[&��W�������dv�oX�²�u����Ʋ^Df8ܣ���Jݑi������(1�E郏�*u�qs�rt��U�34��R�\_ot���s�e��|e�e�#��2�?�a��cd&�k�6����Q�`��]qF�x�M���M�8⽜����D��Ur�"�	J:Tβ��/4�t������u�V���Ǎ��q\۶��F�qa�b��]�[tg<�.@����tv�{\��\qncu��J}��h7=�'�K�!�^���]�5�q���B�nɮn��;�l��Xz9ӯ�{m]g=�d�w0<�F�D팋��덏[��KsV뱶8�f�ݻ'm�+%�3[<�I�����笌�vzF��r�l�[U�nݢ��\�%��ӑ9���ɭ�y��t֜�����!�r�s�PVn�|��x�J�Ц ُ���`7:%��R�t��k,��go&wXx2o���1�±�Ỿ��x|�D�޹���t��}�P��x+f�]�p��. �������K|�w`�x�LEQw��2ӑ-�:ݤF����i9t�9����9,n$����e����`f�<K��;��Z����/}pwH9�(ԑT��e�!��8���S�x��NkxJ�K�ͲgzN$n;�'�i:�L	��K:���pwpwp��j����
]�$��?��ؕ�Y�{VL�
l�!$�^���3�B���W��Iq7�t�|���6"g����Ct�?���'>t�>�$��A���We�l��sy�0�O��?e菉[�VL3]����r�f�m\�iLR�*v��EA-$KxY���A��T�� ��C�_k#>��6�?�F��i_��\W�I.O�G�ӎm�C�Y������5Ybu�:�bX�RG<�c��;�Mt,��G�Я�N�%��Q�'rM}B���*5�ND�A�;�ӹD#�@'�S<��#k>���%��1�f�b�ٍ3vL�]�S���GQ$�nV��Q�.H�6{<ݥ���8�<�x5r��
>�^w�MA�����#�:n�19��N�1��[G.v�Q��!�oe��kr�^\xfq�|�ۗ�lC��#�/ԋ����aѽ�Sp���TUE,�F��~����<ٺ�4�!?^��-|B�L_n(&��n��0�Kp	� ��9����[d_u�I<SX�#�#�s���L f�4��S3)c��JY^��b������? ��I[�O�m�8��=�Zὺ͸��qnn�6�!�օeO$B۝uS&^M�	��,�YA(am�*��s*b���9j�24��+i�?��s��>���=�'>��Z �NPnG�]�w��F$���]�sX3���+�^���L���Ő�{�0c� Y��%q��X���f�����=�����/�~w�"\%%�p��ѳ�ب�u!���^�$�}i@Ӓ�^�V��EXq��0H�
��Eb��dn�Wa�+ϋD�����*Ju�8\+p�)7ܼ>��T����w�F��U�'�ς���/vC�'�t�L�m']]5����ov!d�}�� � 0*�����V��u=*�]�P��ك^��t�=�]Z��T�����TIIY$Q�J"K����3R�{���8�����������#k��Q�,O��U�H����גܒ�c�tB��QJV��_���@'��L���^u#���p5�nz�e�*�QD�2���q�fux����]������r����,��.]xB����Ԇv&�\��e6>J��b�����c#֜#��^��[�v�+����ֈя;��z����6�9�����+��k�:�+wO�eY�Y�Ƈ�X�{�3ɣ7c\���e�^[KkTb�w�;���E�˧0<��u;8ʫ�[ݝTgg�����ak��%�>�N&�`9����a;hWˍ�^+���j���Ԉ��8�e(�m��I+�8�X��-l���s�A�!�SSV�ҝ���0�tĜ9���y��]�2{���	�2Wc�����f�F9Bv�	y���z5�X�w��C�Q��+��c�-oܜ�b�#�d���ށGN ��"yI�][zD�q@�0����n��/]��e5�f8�mӛ�	�rID4�2���p_W�K���)~���~�����a0s��w��YЙR��������;���m�\��l�G�njy�m�nm�z�RyaجU�T��*�2�<�lD�p	�};
�$|�����8���ڻT�6�f����;#kzck(\�=���d�7�.h��~��%�%N��~�곸��W��7ͭ�~�۝��(Q��1dU��g@υ,�Dqs�b;���EɱT��;7q����@�3����v�i���!�&�7=�6E��ׇ�(�&���ڸ�j�����kA��I���]流Ƥ�h!6R";s�^��[����f"�����ًJ��}Ҁ)/n1�{��%�
E�0>w,E%�^��\��2�S79C�u��>|�ɢ��r�Q���Jw6Nc��Sy4�5��̄����7�e����XJ����e�Z&�X�{y�nШ�ژ꣕4P��w;+(�>�9�� vx���dGlU�tf��ˆb���7�����|"2d�5�!�0ᓫ �=�
����yߺ��u�Ľ���A%\ ��an@*�w����
�<��.��D:���z2��{�ӹ~�f��8	��=�ә�${f)��;Q�G��nxyj�+e,�b����:�T��K��2���_}|�;����c��kq���v�=St�S��C�%8,�2�� r���.��q��f3�Y� ����9����]=+9��k�۔������k	e�*�TB�t���V�RUQY�#�¡U�K�U2��ꬦ.�$��Q�Oaq��o�7ea�Z���x@�n-F�v��1n!���s��R�*�&㈛���=�8�Q�1k��7�sp�%G>%'a��.��q��)n�^!�Rf8���=��fMG{t�Oar�gy��j-F�n���{��|�U*N��A+׼q�YKq�o8�|1�Ż���z{���'��Z>�DtDR��L��k�8�!����۫�9��;q��鸻�n-G�RzC�w�Oy12���v�����7�6��E��N�u4c&���`w�ۘ�YKq�w4��!��{F \^ߜ�V/.��w�Z�5�Qq����︺�L��_W��O�J%��qH�r�����|Su҅A}n���k�B��|Ů#P�'�j��D�.z�w�ۈ��Kq�s4�4�$�'{�^MF��^dLR���<�c�N,E�P2���[��H( V��eYU˯;�d&4�&�\{���Pީ1v�̈́|�8�Q��+�����*F���-���K�evӪ�����m����n�	rKR�d�>z��ѪP\
ʸ��.G����qĸ�M��ǏKeB�;.���B�'Ue2�n�*{����uwe��Z���\F�$X�F���e�*�\��h���^�r�Q�L��q;t�w�9��8��˘����E�	��9�e^N���J��OWov��C<�d�%G1�����#��n3XQ�����㲕�+�)%v�IU�sx1z7�P�7�[��#PB�����wR�/"H�t�@�Nj���A<�M�
o��x�s	�*��$�<�����nbe3Z�j�I��Ť���g��ֵ��(U>����1f�B��e�eU�o\�gp^7�����Mu����ZўnͱS�Ȣ���F�ڠꜥڕ�rU�9,��kv�`7�Nw@����W]��s۴w�@���:��q�mRI*j◨���m
H�n�HHK��T��%�Q���Kޖ�T�����ig�.Ѣ�U1Yy����;����tݏ.�/*�Eg��*��o�3�7�_��A��s�멒q#>��.��s�����҆cPp��$��b+����=���Y��n�����Y��Wc�@��v��n�3��}�Z���& \;�LG=����=�ݗ�18�����r%��v��9�6�Ty�t̆1�wt��#���G{t�Z�<��+�9������C��$vQ��*�w�QM��{�Y+���u��Cr(�{t�� �w�[�C�.7ǐ�n���c��hT����j�g5��׮t��L�dT������α {�A�����5��������n%K��2f�b����b�b���G��p��-��Uid�`�:��V�)n��}�� T^j����xc*o�|H�"=��)0��'.J�jC�PuI&F!PK�ؒ߽�@׋I��,��R7�y�M��>ma��u�lȪ��bE�(q�i{�R�J�G;�}%�R
�P�BMLذ�]i!�3X\������(4ݶ���">��HB�
[]�D����E�j	�=�쐘Ȓ����S�'(��D�c��Wq	�5�FcQw�[�cq�sk��Z�D�'�.`�u�(,9�w�p
���$�3@\6���$^g�ۆ�5۵�jq��S�������[���9��$�"����Ut���	frƛHKw��NYm�Uo]��*�@s���}���ߥξ���M�h�F������4��=����*�n=N��j��#)��na���P�v����1�Z�w]�����-+�<�]p�K�}4��o�q�)�������y;�^uE{�R 0�_y6T�k|{��6},�7Y5�Y��_<G��fN�w��������"`m:�+�;;��E�O�6��.C磮-�j�N�΢��Ė�1�pv�����&�I�-���=c'���p@�;s�����T����wF�����v�� ݳɝ�G3�<t��d\ �Br�v}��Z�&6�ngݦ���nwv�5\u���z�x���;n�x�q�9��Z�����%��F"0�����yz�b����Km��ڷ��t5k��k��mIMn{n��6�8贡+��f���`3�rd���9���=�99|���ܶ������6v�{{��M���hk7j��Y`[�����[��y�p3�pv�Ԙ^����L�z0:y]�?pc[䞵�T0����(1q�$s�ޏT��@�+�2p���y��=ë�tF�=���Y�)o��縸H��3���%�H΄=�R��p�g�2������+7egE��W �>x��>�}݉����+��x�8f/<pڣ�s�g�x+�m���[���3�޻D�2�^�Y�s����\;Q�[�iX*l�+u(4�I�B�]<.9���|����cR7���UtuBt����We���\ݪ.�����k��];mrF�jE:�s�j�N���ԼNf�,j��Ri����y�k|��hmE����E���Z�5o��^@�N��{�������)41�Ou��K���j/n��ƨx�I �*9��}�/U����bv�C�h��C@@�#�̽¦����#�(:tE��,���:�c��Ie����#~�ͱ����MdQ��]�n�o6L�8\����f<A�"w{�y�F�I˥���p��]A=�dN,�w�#�vr� q!P���7IQ}�E�Gŉ!�s�Q;�������A!mz	(𵅬r��ImJ��!�d�P$�Ի��{�F�B���}����{�Jk4�}�1���B��e�ؾ�iRH)B�2�5{��|�����׮�����/	�!$�U��t��B���1	�5Ԥ�)*/#PK�C>A��H�ϵ��1|�7�HM
�/i�#��z}��-�CQ���9b�*ߝR�J�/P��(h������D1�؍n�! ����1�7K���Y�y�{{.^@��b��	Z�����xr��S�S�����"3uWl3�� |�b����wXG�O@��#�i3o_b��5��B�j�d���LQsH��ۣ�Pwjp������TC^���G��1D� �u7fQ���c�GP>ﻛ1�8�=�7�G؅�|�#��r� ��S�C�}���,ά��v�Ws�31+=؜��Ѧk�'%�޶�������D>,]�ޜ��s��9|�ښ�m�\d��t=g�����C-���!K:�)-P�),�7�aa����<ɑ�[�qB��
�r^R�	V�ҬU}���1�.�`t=���d��~�e`8�.�<�w����gգ~�K��KMT�3 �R�Z�#���t�%R����v�$MDB"
P`3^�����/�7_�����Y�4�n���0�gay����ȣ��Y��@։���[���c�����+�����#�C,��y��y�O^�DuK����%��%�V��(氟`9�F���q@�wGr���0�>�?*� Y����zșF26�h��3/W����{��y���@��2"�2l�Ƙ��Fj��W��޽�a���H}��d����69l����[�ֻ�L-����0��;�{����O;�t隮gk�����q����w��@	$����i�_y��K$m�dQ�Z [",pr?���Z�]3�U��Ǆ�����L�Z,u8�#��.�'iG{���V����ب�p9O=�t?K�)�DRm0KZ*v��z�v����뷷`۴.<�r��a[S������b:.2u�4�CD�<;߃���R@��%@6�7{C#�;�쉸�D�!�/�>��sx2�l
&T�\�s����ʽ[g`F��crǯYˌz�nr:��EN���S]�7�u�k��lS��vZ�t&>�M���C��k����Y�I��2)"w����u���ȶUj��;�{������Jj�����r�Zdi��%���r�ti]D�']�{���q/��]�7�\���!�N�FF���q(d������1��{�/�_t�q!�S��t]n�B�ˣ��V��C$�w�$�U�o����H��x}������Z����:�=���`��k'=a�(���G2�r��]�8��'����w?+$��p?	��ʱ�O�]"3�ӻ4'u:]���õ\�}ں��M����g�+QEh��qw .��y�㍺�Y��g�b�<�)Ի�Y�s��k)��ͧT}�{p,T�n܊�[a7�0�\M���yk����Q��r�ĥ����s7&���J� 5��Y�A���^�b�jË�t͸3Zw�h��f��a��c��0�������q��g�G*�z�%o,��8h�q�=��|��;��\���{��P#mkַT/2�B�[�G`3["؏�OaPw�=�'=�k�כ�
�rj����={�����(!K �Ej%m��1��O��a���@���e���F�#WG��t�w��N^iE8�<N��ج�ɕ�o6�:/;��}�xxF��������!�k�4@�nU�X7f Me�y��6�Zw��\-�(���wｓ]X�n����-��+%֊�Ѱz}����*�oCS�z)z(��f�ͫ]a�l��q\�.E�a�v�%�M�6��[�uӷV�(ꗍ;�rG$�.�UU�*AH+
Bn�w�;>���٧-�u4��c$��V�{�O���ۦ�H�����Hy<<�4�%n����\�e�֣��=���W��r�a��E��f+��,��P,x���{���[��u��΢wGrp6�(�"��U�~y�Z"�BA7��Ƿ�޳�/˝����&L�he���i�k	��Ǩ	[������|��eȤ����N)�+�x�1�`F�V ��0��F����{�tg�~J�/.��G�#w]�H�"\���kU^��[�O���n_��[*�8瀩|p���P�� 0�<ݵ�)	%v�	H��2-,3'���A���B��׏���ڡ՜��/⟣J� ̀x�\����gg��*qZ.�LL]u��Mp�د � ��A�@�������v�O8]��6�j"�m�E��
�Q�~>L��;�{�$x�;�TW�?������^�녑z�2͏�qHq�Z����,3�)=6u�o�#sD���;1�̇\�_6'6ue�.%�eo8����U�������t�U���ذm�[mU���[o&w�`�Bn�%��Imndj�Q��_wc��ww7�e��v�q]a,�خ����l���|w�xb���W��M_�í��~�οyf�R�k<�K�L��0�i�VՍ��S�y���t��	߾��"��Ͼ�s9upj)��{���@�e&Ux�����yμ���qy��'W��2q�>}WAF���V�[k�z��B�v�9]V��UQ[R��{+ӕV�n�h�;���[ϒ�}c{�����u��1R�d�]u�d����-{����m��*s�L:�Zڛ��H忦��,�e�+��j��Ĕ���N��7��#lq���Y*a<pu
�{�T�Q��Z����<7��ql㽕��>&K��Kv��*�����ʮ��Q���[@��s~]N��וk��}�u�}~9~{^�n\Κ�R<F�w=�y(h��s|�
��rVSe��PMJn.q	N{��C����d���A��VGx������\<�@���xb��W��v�V�X�#�PA����҈P3���h*
q�(��z�
�?x��7��j>��'����Sx��h%�n�f�z��ѿNf1tg�߻0�/�\���Y�W�͋m�Vv�q�zF{��uf��of�FP���M��H��䴱��,�cl�۬'�#ɞ�:NR{�L�gb3�.e���f�Kяhz�E��F��茂���u��j1���w.	�DS������|���0�r������f2t���d��ePU�J
�Pjm#S��<yճ�u>�-ÞѶu��<ώ�)o<��Gn,f�T���x�ݥzy�����q���8R�����Z��ޭ�s`7O�[wbb�6� (9R��E��HJW�tMq��̞�帶�kl������q���ahMVp*(��a5ۍ�aQ�{8�xٍ�<�6ܩ�5�fz��X!8c�ѥ�]�;�ù�x�5ۇ�:x�gG�a7+!��q�j���IU�c@�m�Z�9n:�MWEk�#6Y��wU]���ж@��Zn�{��q"�����*r��r������M���_���oC�W��|=㒧�9�kF��R��#|u-�� �3���y}d���2jor����ĸ	w���k��gv��4w'or��<���ܺ�;Y^�p�ְq�Zբ�����颰���ֳ���zy�$��SOI�����
�BP�ӍP�nuZ�,�Y��:���^�\k]:�t��[�]s�(�gv�ALT�µ;�=�:���9��`�o�8�mdSu���-лa�h���s�L�]Rg����q��!���7�ݭ-�'G�����Y��1p����$x��UZE�L��e����G]����l �hQ�>M|���پ��۰��C��A2�+���<��N����+�{�S�pټh9������=\��������;��A@�s�v��X��p�ďu�_��VmZ'ʏ}W��1�x���ϊ���{v�mTY�j��v� ��B7eUM�wZ�����{dZބ�|r=.�:�^F���}*����j��k��k1���+�[е|��	ɍT�o��}%�z��}c�]U?�-��ED��`����y���!��]�`Yz�{�5����Toś2�hf+±�R��yf�9���:F`{�MhSW[fz��3]r� H�11 �

;�k\n�P�`��x�5�/���ය6�R�Ge��˒�UR����U?c���<��TiC>�ˎ��鳦ܮͪK|��%�\Y��x��$>�����0**s��\5��T�߮��L ���EEF�H� n��,w[g�6Y��E�{��C庺8�k�G���j�Wz]V�ۯǯ���0^;���"�9��Ͷ�f�Fڒ ����~kV{���-����LF�N��7�g�[�\h YSa�Ɍ�o;������
��v�/~=�_��M�D4���ks&��PD\#1��Z�c�f�[˴�9���@Q^�����/5��a��;0ç�	3���^4;�h�^ڎ��-��ٕ���mdRZ�E�+d-d���У/���͸���v����m�MqP�t��lДt�R��uf�BwU}��Q�6���,t��4	���7o�t2�|9x���S�P�b�+�ut�mK �e�:��`E"���:s��_Y���xR���~��sz�i]�Q�N��~4t��b�7�pGd�SF�!󿫁�$��0ƙ�k�|G� 	l}����cZ�x�f��lU�Сbh�KpY |̈Y5����{�-��p�������U�G��33��M�v��W����:T���x��G�9��1p�Pc�v��b�c�{��Oc������gf6Uۑ�m��6��v�η�%xHA�.n�a�1�1�7Ov�]�Wh�S�j�l�}��wcݏx<-��n8�qA��A�}�:�ꯣqM�
LZ ((�r�����oc�Y�^2V�4Б�I�����C.4� +Nc��oY���Z��8[��Ÿ�{�}������>z ���%�īkp�.���@���F�߂�3���;1�A}�~M޿rP3_�f6���ȪW�}Drxv29b��R���L��E���d|󉨡����w>n ��)/j�ݛ�Th�J�+�jZ����8���������������*�5��� ���{�}}�#4)_E�>�a(H{V�0�^�^�o^ֶ.��L�ם{�u6�֑�X�}v�~�Ջ|�.��w��ȧ��ލ픱X�t���=5Byoc�\]�޹��߷�N��M�J~񶸒�=���b������m*s�<�J��]��gc&p`�F�[T*�Yq�2����F���rt����띷wb�}�Sd�a��k���^�?t��E߻�G{-��Y�V}��yN��!=Њ�t��
�K����f�Z�I��n����I��}MO�O
�ͣcSzi�N�K�ᓯT����4��'n]��{G`��t1�=��~���o%}~���Dt�{�~rq�}�[��>���̫�4��x��Q�sK�q�O��H�bZp�=�ם�ˇ9��U��)�)/�/��u�!��~�W�Gr��a�Q9��܎'Ue"Tj�,�m�-ia����C[�\�싥3z<�����w�L�vDFQ�yk���$�Q�����9�l�V(M�bؠ�$x}L�U�5-�MLMIۏ�>a'])@!P�RC���G�s�(<a��e��7����B}�t�\<�<nz�㮩��(�]�M3ˢ����;�m���eL��]����QQݹ;<�i����9J�i�\s���91��֧�tt�r7h$mB;�K�e*1�PUZ{niT�0�ǊTʜ��^���0�{L�Z�>����9}"�I�=w�)��ϛ�N�3�@��ˠ��6֣F��{j��Q�^),N'*5 -��o`�w|$K��ٲ){s+,��˔���j�0S�ܫݧ|�He2�%h����{���u��i�2�u�|�0ö'{�q��]��cw��c��B�V[(8�N2�/XNP�	��C.4�:E�kUyO�Ra�t�����U{t�������%AUw����X�C󔅗�K�>�h�Ľ���XB��A���Q2;���ǎ��3�p�v��q����=je_ ��-4����K��3r�toL����q�lF�K�	'�h
Ef��;��k�ұw��X�d��M��1j �siM�ۑ���Ϙys���d�=h-�DX"ȉ��M�^�rP�qO�m�|d	CJ�����1�>��q�On���kھ���0��WBT'(藎;:���nΈ&���{��傱�1��Z�Gf�v�\�=������ps� @�� �S��{n�i�ԧn8�E��,��٭5�K���, ���P<8�>��$��S��x1Ma�kۼh8�.H��^��&�"$U
�H:���K%E�L�ma��l�s�3Q5��a�� �,�FA����w�=�v�D$d �1�=;U��={yƹ|h[�{+���k�ҳ��<�b�#p|�����>�r�$��tr[-+R��#��u���CHˏ+ǫHV���=7�(��s�I��;sV�b���۰ij������}���LLH*�Tm���,��d��0�}���H��]qP��XlZ��X�ʴ��6�x�jwޒ_kxS{~�G���Y�F�[��ͼ�&��ug�3r.��Kˣݧw��x�	��v� njo��}�`!T(3s>�⹏,��M���ş!}��kvB�
�9@dK{�P�����'5�]��d|5�oI�9�/���q��/ƍ��[��s�-��S?���_������@ P@�֠*���4�~O��eJ���P��a��-�xZ �. � (H�   ���H��?�T�6�
 � "��@d;Ĵ�1Rn�(#� kQ���1�28eD�TH��EJ�
��B ��B� !��"��H����UT�q��*H$@�Ԑ�(Z`Ā��ȁ$���j�H��2"H<�����v>�/4'O��2ET	'O�s�Uk?�?o��G����ߏ��J����ݧ��5�����
1߶�8>���

�|_����|�}?���*��T��Z���c��}���L�����O���D~����1ߺ~�O�@�������N�͆�"�b����"�ۑ��T��� �s�o�#���p�AL�E�9���`��"(H! �+" H����H
� *�""�)"�(	 ���(�((H ,��"�"�  H2!"# � Ȥ�"�H?{Z��H�$��"2�"�"�I!�
�$P$dn��KG��忲�����?��?tA@��Јů�>������? ���'㟼>��>��G�/�A�@U�AO������@�_�#���O��X�2��?W���'ؗ����'��|���?���}����͟C��XQ�_���?�~���i�UC��@U�A�?b10���"}t8��#������G�_���QH����:P���U@�������g,�R���>t����A�\@�G��~@����?j�����~���k������>3�8��(~��}�����>�!������}�-@Ux#�F@?��?��DP>a��r?�͞l��8ؐG�(
nY9��޿�u���g�	�?���ɽ
�_�=��8���n��!c�G�k���O�3SC�=��^P?���|D����4?��C�/�Dl��sJ�Y�p"6}������-���k�v����_��6��]��BBc�e`