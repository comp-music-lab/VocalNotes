BZh91AY&SY*���_�px����� ���� � � X `b$�{�    =         h��      
   �            |                                      ��U  P  �E
 ���JU*�J   �H��%@ E  D R�J  (H �       zS�B�ۀ���\������<���X��x�� #�=�盩�way�y�T<��t #��������㡀�T(�Tm�>�S�P��r�ҔU���d�)J���O��>6�xގ��*W�\��5ޞ #�J��^��=�)�+��:���/���B�_|���
D�       .rB�����R�,�����)�'��S�ҕ��t�5=k ��U�n7�RU�<f��iJ�����ԥ*�����
U�^/sRU�5=�"H�UI,� U��S�iT�5rԥUϯ ��R�LM�R�M/�}�J�3x>�����R�� #�%FZ��8��4�<�ye�S>�^��+�@��UH��       �5m��>z���Mϯ�zU>-/}_�_-J���]J���� >��*�O��5��������{�k���yp ��R�->��R�������
)� h�I�{U|�U|}�޾6�����A��qy1���� �F�LA�X9z�ZS��w�ҟU �J�P7       t t���8=1޳���;�����}� ���̰{4�mm\ZQ�ۼƁ�Ѽ��z��/1��QB%��@��=Q�9j� tn�Y��bת�cͪ��rP`у���^���=���Cӈ���)�[�      �JM��p �3�2ХV-Q���
.��W� ���f�s\ڡ��x�1��mP <N� �X�>R���� DCl������&� q;�m>���_6��g^!�V`h ��ů����4:�����T���      @j���R��0L� �``E?&R�@И @0  ��4�a	2�T�F�	��012A��D�*�	���     ��'�QB�@@   L��MT�T����<���� #hd�Ї����~�����|��5��}�r��}�s<�?0 �N/�� �I$�$H~�H$��?� �I�?�?g�,�� $�?��V�o����[Um���ݶ����H?����?J��~F/�`��i�G����J/��5��s�����D���&�&�n���t.%ZssN��v��Y�i�y�+N򢞿=L�R�ه9-u��j�&�T���n]� �y^�x���"Q��ol�:�Ŭ�m��3(}�1B���{f�nH~�Qˆ�{7�R��xNSr�;FG֎���EwGd�������t�q�R��z]�g?$�lY�������%��Xא}e"❝�8�n��j}G[
Pf�ɸ����7���1�7')$�P�J��X��%�N>+q�Ή��Nίy�_c颦�㴮�۔�nu:����L�4 #Қ#F��#��:���˺Ma��q<ьG���|��]핓��5܀����w�����6jf>�ٿ.ދZ
]�&�v3Cz.B��R���;&$$Yͼ8�V���9٥e�;ND{5s���w��ܹ��h��#�������&�׈�2�y�)4��%{��P$w�Wg.GH$v��/	���t��7L!wn��&����#.�KcZ���go��G����n)��WO���y������k�١d�;vn'�������q-\����d�ڷ���ǡ�g:wz���#������>�P3�4#����i�Xvi:�cGX;t�"b*C����(9���HH�Biu���^9�^��2��ZS��c=q]x����nh���+9Y�ἚCf�oǀ7ou���]��ho��3�=�뽵n�;L�C2��/�3�(�Nu^�b��n�n���,����Ppȝ�Uĩ\F���k�c�!Y0k��z�ٯ;bɔ����Dd��KTV �۴�LN��+��"�)t�u�t+^��X!�(Ufϖ��.{���h5V����G���VJ�)
H(�Q��Z-^���/I|_W�r�ٹ����⽝�5�B��{X���H��2�E���c7���bN�ӱ�ю)ho MOMA���؜�B��mN��]�.���G������̱[���S{SHV1�����ӛy�^Ś��� ��/�o�!�
t���;/���`..B�Ua��xM�b94�%�\׭]�D����e�cЀ�]���M���S�M�+��(7��v���=T90Er�2´���8�LgJ+De���X�	K48F<\T���nl��ww+Rܝ>|u��.��ly$��H�t� ���<ŽB��b1jZ�{�o��1�ScN9����5�H+g&�Id�@�,��P}hx���툽.�%bCv�.Z��A�5�/2`�YI8�&��,Ȑ��bq��hm���՝�l��{�叝B��Y��Z֐N��W�~�6��۝��)@Fst�2�	�&���Ӊ?=Z�)Xх ����P�s|��iyʮN!�8��f���7�gn���w�]w�r�m: hrս��\n��v���'���B3t��_,�S �����o^/p��q����]�k[�����E]�� n���1�\\m.) ���`����"��n#j�	)�F=�v��h�V\۝S\�pO����*|�����t�>�y�0��虽p�Od��漛E�I^Le�h�짢vH{Ddd��ei�wo\�A����>�ڈ�^�a��3�2o�͇�9���q=\��XkCm����åhE�;F3�D���U�|��n����m9YxE�e�C��d��]��Jx�c�U�vgF4K��$�aWu�i���gG�R�X�����W�L�U��=�n�U@#����=;;]0scUR���Z4�Lt`�l]F�8��uos�md̹N���n���6ePp���ӫn)��0m���p}�6��lG6���X�v;N��:yw=�A�(��kb�q^�F�(<q����ǹi�H�o���פ}�Gbu񓹱u���|�AN�'.ȥO�2�i�.�'`�M �ɋ;a�%3�����dӐ�*\�l�9��F��1�eÆ<�����z'OG�t��@��8Q�{KҦl���V�����7qI�g�
 �ȳ��qQK��݂n�*G��
=��+w9�8�V�+4E�۝�D�KDm�D^���^�1���L���+��]l3�>H��ۼإv��y�Y�	�� G2$�X���|�zSJ%y�{�w6<�+=��S4٢��t|�:��һ�Nv+I��u�1t4PA4oK��3�J5� -�[].��O�d�oL�r=��:��w�kƛ�'5�M��Ø$V�U��ή�fG��7�ߞ	�N���7�c�[��LG'�3.ef���h������fŠ��+��e�Y�B�L�7�b`,ζ�b#�x�g#2w*W�S�g;�m|�>{��q؁�q�0�v��2�'gij�a\N���5(K��@�=�S;�˝�V�D�˴QA������r�6���!�wGN#��c1�	,���ʺ�\�{�PL�ǌj�	��bK�vI,u���	�s��r{w�$�IF��1wj84�E��U�M@!�&�ȶ��cQy��,J�\Rk���y��'#���BػM޿l�DX��=���^\�x�W(�9E� ��ݽŕb������C]����+��y����٬'ưp`���.��c�+@�6�+�p�80C���:\�4�F\��N��w
�pO��!�?����㥹����@�u���{R�ݼ~��[�]�M���ͭ�q��&�Y�@T�.mM��Hu�]�:���콍(ӽ�^�7ZZ[�����n�u��.�z�`��-)�%I:Ǝ@���iw���]�R80���v�;=�lG�QF�x�f�xP"u�lA3*y^��DƷ#ǫo�.v�漽��w4�4f���L�����۝^8���� �����p��v��n�����4%)��B-��Q�F��㩷vE�#����ݽ˻K�|��5:�a%�R{��"d���r��rX�8��-�k�չ�W�t�<P���c�VH��y0jd���(hZ׼���cAN��L4��1�uA��y]6�>�5ԗN���-7��7�>wb��U����6R��5�J��,�xm���rm��&	��O#�	}˛�J����D�00�"@Z�ia���b����I�����
�p�w���lw�
���r��p�\���6#��lU����5���������n�psbb��H�i|�c�M�>�^�ŕ��8Yw6��1V�����7ooc�:�}�A�n�N��X�ELե@�|MڨZ���0S6�:�	�w���o <U���Z'S\2U���ok�f��+|��X<F��7ypf��V�>���n3B�vE��ط4����Z0:�[�2f�; ܛ����o&�p���=���.�
���S5�M��ٺO#�V�9JG<Q]��óz�a�;�ٸj�p9n��+�;��Ӄ���v�n�#�L���O1юׇ^K��(y�Ǡ�ivo��9$gR�ON�0t���H�ãWZ�^�8�w,��h�3��k��Z��p�xk�&~Ի�Gy�{/|��zm �㘢�e��m]X2ntl�ۻU�X�opi���xt�{x�:��5n�L��E#��W���pU8*Ʈ����*T��2^ȍ!(Yh��o��I�˹�jx^<8xL-�9�{No>��1�o/��F���R��$�uŔ�:_e�Q�uI��U�s-�f���%�xT�=x��r�=,��-˝����oZ�mٝ*r�T�|X�5v�ީw�����\�f�y���G_�l9����^�l���c�#��s���Z�wD�3U6;N��{����˲Ɩ/U�0�f@˸5s�-�׶���	l�A��|�_n�h6��	�5B������f�J�� rŕvQ�lO���:���1�����L�f�7s�eU4r�o����wA�z�o���u�g-=3��5�p�u�+�-�j�>���R�}�ٝI�q��Y;"S�0bP��/XŖ.�
�AQ_vwp͙�=�vu�d��ER�pD�t`j��D�8�E�~x8M�Ћ���.ӵP81�=*)�լ��l>G�׿3@��^a�MK ����������]�s}�0G��i��&��=d��Etۄ��y�z�Wf�*�B��u���d��J4LŽ��k���Ӌp?��b8z��������D�v��CI�R���쵭rگ�o P��B\vf�Ś����\��WZp�s5�WMdi�{ ��ј����v�h��m�\�t��M��m�坝ץY�Tҳih�����żY=ݕ�u]�0@�Ν�n��h�'>��Y�b&��#�T��،�ƍƗ`i��3�F̯�T^!�S��;��s}�b�|E=C��w�c n����<oF�yC��35]9�#Rɧdڱ����VZ���7�lGQ25lJL�[�,z���3"�9N�>7���x�
AӨoׇww(�k;�+���6T���b��1�^����9MƗr�����Wp�V��Ǘt�dE�|X��lۍ�y�-�������`3Dj�}V<���q�A!|&>��/N)����Vnm���X�}����I�܇�����nX7w
��*�1�	M.�Q�5u�1g88��1t�:6R�|�j�v>\��4���摄�C$�����i�5�&AS�&奎L����A��{��|!�ms�o\�ePѷ�.B�oC�v���C�sy�ͣ��nuk![��Yl�w�B�uCn��^m�~��D�d[״�ы+��K7�\����R��;�����eF���t�N�&tZ_s�³�}J�1ٽ�l�>�c"\I�|�"m	�zѹ��2��`]p<$���J�Xx�{"�N�,콪�9����kxd��!ۛ�5Î[���t�M�{�|f�n����\�k-��'X܇�iɛ�\ۻ�O\\q<j�N�����D�Dj][��y:���ʚr�j�T�:]�M�u���p��c^pV�"k�vr��u[���\� �V�S��u��%�hZZuV�R�*RXӧ#ٍ�]�5u-\@��LS���ܒ���syzYf�pl��d˚r�A�
��Lj��V⢝ޛ�����/��Z�B������I�d��\G�"m�˳yS���2��y&�o0�Ү�鐡�D�s��*��%x�&��:u�:r���g�����B�����3O0w���Q�}��t�����G����(�w
x-Y0�	��:�b����կoM�]�M%.}��-7��hЮ���;���ND����"'v��j���Y��T�E����^���r��Y�9G�潪�L�B��_
��ִ�n��%;��'k'���n��/Rp��hR��9��l}ږ��� I��^�>;�6Y3a�2n��Aծ�Vp|���_J���|ȅ��/Z�e؉u�6r�7{]C�����Ի�g���"7X��,o[Z;�f.2�̸U9ok
�GwOeG�-��4���T��q�ykVok��VH�m��x���c�V:�jI{��K5��\�,L�)B�KiW{3sp%��W.���#&`��Z@~5(���Z�Kx���"�����+��3���O6$�#nj�ϳx[mc��c�1e��D��{�{�P�Rde�xoh=�� ,s4�ۜ_k�0$Hz9������=ۺhdsd���o�@�K�U�e�����@�}M��ћ.��@������#|Fj��������F,�Q�K6���\G@���b���Z8�f�U�e{3Fy���y8e�l��Mg����66)8 ��V�ZN�X�{���jv��{�>��	��爆.*0%ȸ@՜�������౨�LeW��ڷ.��ٽ�K�5�Q5+�g=���x�٫�PyV���w*bM�{��Z�|����kk���Z��M�u�Yw[}F�ݙ�'۬;U]P���a��k	���z6ݡ��6a�l^˄�U0�0x�l��67Z8��7q��Y��8��XZ� r�aĘw8��MX:$w��u�_W��n�c/��]+�[�=ڸ��m�-��9��gS�d;�29��u�ӆ�Y�2��8���X{c�>�h������*n���`׆3Q�l�:Dd�a�NO�N>�f���7�`!ߎ�L��a	�U�<d۵�`�Em���^��-!سh��a�z.��Q�ͧ51�#��{Ӌ�v
�m�ۣu�6�t
op<�N�JM�	f��0��b�T�i�H�3p���a:����oT��nu�Vk���oF��+��aQ��i�Fn�7�۷V�(���t-��hAl�H�cz�Nʈe��>����i��a�e��w"+q�8��-2��K���YvP+iD]�\�l�9�]\��3Or��K�y�<zv��d�A���O*�:f��g1��$�va�ڎ�;7�T�t/�6vZ�Z��5
���x�i���'�!ף18x��k�3���Z�$In���"���%�N��ݻ����^�� ��2,a� Ҋ@�0+�k�B�!��������L�A2�S����=���*���O����!���x�yΩA���z��n�U��Yk��D�c�Q���a,��
I�ʱ�`-��p	:�;D�N\�˺�%4$O�n������]�+
�s��]3�%�N�4���כ5��i4�0��w7 	��r�AO�X��1��}~���Ubj1�����o�R?���b?�(�Z$r��ۑ��d�rv�n3�H��{V�np�u��m9v����n��ײz�s�W�����-���]FF���������n�<�\�Vw=����ã�ll8tx
ڞ����rarZ;]�ۧ�\v��q���#���t��^���ӂ�-&:%�0l��m�n����2dE��݅C[X�;:
�>���ݸ�y�9g(xi4:���KJ�t˓k��].{d��J��d�������]����/lv�DaZ셸bc\�����)̈́��keו˳�rE������X��N�q��y���%�Kѻfǌ�ں=�m�U�;p���[��z���srf45Zva�m�5��렄66����>2Wn�c�.wv�vł���bLg�jqS����vumrvJ���5�w9��oem#�ݠw�����';�]���lN��Mќνu0���v�d6���k�v1�\C���;v���A��m�N��B�ܣگR�ǭZ@��.�/�g)�iں�܉b�OW/��v��]�2�s�p�z�vn�c�n�J85�aC��.�T���q&�8��f]���<�#��<ۇj���jP�᳼c�]��L��Q��n͂{k���96N�pq�^wn<��I��FC�y{70�iʼkc������v��D=�3���|{mNϫ�mv�;]� ��5�q�϶�㥶%x5�u�k�ϭf�N۸�ӫ�N�`��˖њ�Y-��g2�����:lc�g��]��<!���mpmWr���lu��	��X�%��P���N��㳇u(pڊ���LZzM6�]�n�~��۳��q]hv'\=������\���'-1˶���6ջ�{<��s�d�:Dy�����������7.�ns�ӂ�gf���l�: �{'\��v�z�,�����269��Q1k����A�[<��Nn�J�pXv�}��kRlh{<Że�������c[O
����ۜ��;q����Y�nP�(v: 3NǬՈ̹Kz������`���SW-�;�m��[�PE:;I�=<�Ѻ;D�=��=�P�a�&�"Nk�R�;{y�o} ��$']n��������c�!arN�c�[U��wl�#�:6y�Q֞â�7;n�nzL綰J�u��v���.��6H�<6r�03�T�g=�zvkʰO�^�7и�C���|w&��7v&ݵ�T���+��c7K��x��r	�g�aɶλg�Fݘ�`0"��)���ݺ��x�b^݈f��:�rQ��d5�󳭆����<t$e]ŵh\�<v엫66�����r+\���9�]|s�|�z��֒wa�9M�}�_3�=�._8۬�{-��m�rtg��K�ɂnl�E�]���`K���j�y6���u��[WX�9ٷc�8�K��g(X�8���V��0T��{qn����sk6׵�n��vS��v{�ɮ0�0�=�l�bE��N�[����%hSu�t�:v��b���A��5�ٮ�b����[������ٴmn����li��\kN�9��l�Xз����<ɟ'f۷Go�۫�0�3��:�J۳s���[�+�<�`$��kZ�Γ�ր�pM������s[v����_|h��HmCΖ��wKV���#p���ɘ�DSһ�/j+FFSh��D5�էjۈ��d.w�5�{u��q��GK��*U1g��U��;m�Y�H��n&��L�l��<��0ä���<E[�!׍j��ԧn��G��&Cy�us�������-��3p٫pgF�Y�L���'X�ך.��f�[��";b�s�gpuv�����hF-=s���筗�T�w=��<��u��3�׶	|��\�5�l��g�meҰ����c�4�.�I"�i�F4t�����q��⋁�^ێ�Ӣ�;<�[}}�;���؁ӝڅ�����a��n:�y�2WWn�`.9������0�;�,W/m�n�󋜞LK^n9���k:r��3<��ڵ�����x�8h�̀h�0u�lh���l����;<�ݭ��!�x��fMМ���>�����V��Q�nD�987n<ݹ஻��� �<u��`����A�u��nޥܕd�V��z�v��sh��U����n-���j����Zo=m��=��\���u�`�m6h�i�������m�/6ƶ;Aζ94��';�L�m̻����:�üa�f�Ψ��UG�2�9�7 �or�;=��cv��tFfBz=Y��.����͂�5¼�R�v�Ś���gqѤ����q�s-��ݭ�u��9�K�G<\��l\��ӽ�.�=���rh��q\�`����$��X��>�a�s�v�ݛ<���cu��3�:��m���T:q�홥�=O`�
��T�'i\2�<���q�k� ��;bOl`�h�
���g�	Z�v�@tCz7U�� sj�q��`���)"`�\���]��^��v#�k�q�8b�C�\;��㎳u�����Xz�zx2狳��۶U�mٯZ7!���*.v���q�p�7�*-o4m����Ef��r鉇��6���G�n0+�Z�P�O88M���m\o�_q�}��aӸ�0d{�ծ��йlN����@Άs͘�X��;�A���\�/v�6��}���5�e���wm�]����k�\�=��sЃ/+ȭ/�.m�^��3ӽN���kQ.�<�s9�O8�v{P�Ƣ��h��nН��;gv�	�������k���&1�-|."��=�gf�a���nYۓ>��z$��0�Zz�8�#���vۣ���6�ݲ���q��9��Qԭl'&���\ݲ��<=�ʏ���ʤN�X�ph�ls�j��UW�	�8���w�%y��m\���q8�x�쭗N�m�}y���p�/N>l�6�C%�)�n�gVC��7u��z|�n:��<2����F�G �������p��d��F/h�q̝qv��G<�nn5ۋ��z�zv�*�6�]so����N�ݸ�Q��N�ݵ������������Ț�;�7m��H\v���$�gGc�=f��]�{%�6�u��p�c�<���z��'V��g��H4&�v�� ���q�[�n�ۻ�3q�n���۳�٢��&���f��局�3�m��s�5�r㳶cY9�A����/"lJ�oI6�FƝXyϬ l�]�/Z��6v�8:�`�n^:w-�u��z�g�'V�٫��xK3٫r��Oa8K�m�0g�.��F^"�y�'a7ok��k��!��]�^;j�n���݇B뭝Ѭ�'ek��Ϥ��)�1m���y�:�;Nń+����}#�d�;c�t�Y�Vv:e�����-O;vz�K��6�7vz�b��zq�v[z�F��h�o=v�m���-���M�r�n�>`^=v�����6�n=c�뫮����|��6y�yύ8�m��=���{[[lA\n+�۳�n��l-�ȣ��vك��띊g�!\t���ch�%g�R6ɻ;n8���65v~n���������i��#���n�;.��bg�5^�}N��:,&x�N�f�<��i^�4o;=�qK��Z�<7l!������[��]s;��Q����b��wo��Om$nG���b���)�m���\��qmm�����g!aԼ����6l����T�P�kټ\{nK�]��)uv�`�ۃ(��3�sܮ띺��r,���6�.��q�ے�9��̛sA�i�ܼu��^w��x�Dny��`#]��ln1O[[ue�B�k7c`��AT��Y�\�̱��(�DWB��F,VA�	k÷]%�3��dr�����],�<Uа5���H��Ϝ��ݸ�K�lɟ]0a:N�9�z
��s���M��6�]��v����0���=�=+,=��>K���E\k����KG'F��f���%��4:72Xz��\���6��q��۪8ڷ#��:�;a6����v�C�t�"��gX�p�qV��e��m�M0��m��¹��Я9\��]�h3t@��|n�����:[�nNy1Wv=��/H�����P㸎���n�������+�յۛ��/i�lnw���t�v�z�v�uq�=�)�8���I��=�E�uqo����-�0=�F�0ub�֞��Ț3mI��cCo[6���<oB�cn�6ݮn�lj�vp�s�\��x���y��k!��/���7d�iwq���ۢ8���_;w�n��[�$s�+�<���km���^a�QC�ݪ�ېn�f����\��^��v���y����/Hݷ$n���pq� a���8���֮9q��à{�����n� �7��Y�,󞀻h���A�٭��.�Z����Һc4V탵رm��{a�s�ܵg���e�!�	�F�k���2[&���˼.ۊ��s���cC�Y�#�m����s�4��χ��#�8�l��͂��젚�3��=��@��b9��=�㞥�.G��#�rD���Jkt�pٟ[4[A�Ys�#`9�������h�ݭ�L����=s�G����l��g�E1��]v33�z݂��y�Jz�ցG��z�q��o������>L�x�v:s���۳��7.۞À�����O�u�N�j��gF܏o\�����+������cK�rv\n�2vx��k�ɋH;\y��	ը����ŋ��j����wn.]hU������gi��F;n�ϡ���Dm���	y�j[�<o��	���I�t�pa
m��&"ܦ_�۞�WJ�9#ҍ����*7����]7]ZM��V�UA��#��O៏���A".{+��U�ד�V�9mȝ�Z�p���pn�F8w���;��7:��<�pY���/sr���t�u�-�n���9�uC6�8-��s`�<sq��^6���6�2�:٬i�#�<�=`�P��a�6��۵cv��]�t��V���=���;������FOV�5���K���]\ܭ�#LE�/s뫰q�����읻Y���[;&���ɑ��1��[]H�nv�A�����)@p0���N�.i��>\��sa,b@}a�y��v�V��1�t$����L������ı����~?���r�fd1w�{�U�0�K���z�A{�fz�"���$kJ���v�&����X�ZV���jj�,^��z ���9��[�c�[���q��fȉZ���u�"�Sձ'�������>${J�l�pŽo�����0�E��F�kf��:ܻ�E߹��?U��;޾�М�h�t9���\$�e���>�;���	�Nk.���Bow�3��`*m�2�8z�;��-J����%\���/1^�&z{��1�Q�p��`���
|`y-���kh�[��0voP:DN�t=��~��)`�����8^�}@uiޠɧ㢪w�^��.�_���%z�vj���B+�2���Yws���O�㱓h�>.��~'��z����.^^��4;݆ALow���--i�|��zpOrKӫ��k�Gk��D�|	y�o�w�{{n��nvP�+���n�-۰�ѫ�	��V��%ú�u�D���E�F��a���^^8�3+7{9ΟHgn�:p�U	��un.��"�>|}������������ڍ"�wa���K��Q�&謹�\]�m����炙9e��#V������vB���,W���,*)ug�X��W���6������������k�|5�L�ˏ�_/? 	g���C�0���#����q��Noy��/�Ia�qO�~1��X���N����z��϶x=:��폟���^�6tO��)Zq��8{�f�u�wU�j��̓���d�D�)���\�׻���(;�Ò\^�<��}5d���P������o{u{���Җ��Oz��<E���i�X����:l5{K��8�~���la�����Ezz8��W�?osﳯ�,N� Ӿ�ú؝B���7����t#$��?{��7��/Nǭ�I�B��d��ށe�+�zQ�)�;G�>*H��T>����g`��㎘Pʥ�X�A��$,��Vx�z�&���u�?�ԇq�B�w��e�ky�,e�͈��w-^O΋2�^��������z.��8S�Tk�6!���Vm��V�	N��}�Ƿ�6c%Q���|p��Л﷾��N������	�<��ȟ�ۋ�J�ޭ���~���>Lk����������hS�+���Fjۮ.�h��.�(�\�}��V�w+^����^�y�m�>�>Y������wnY0`�b^h �{P[�V�\U����sy[(��zA���z���ݏ3e�v���jcS�)����q����Q~�0�S��_z�7�{��ŭ�7}�()�lY.����k`�T��ܜ#�,�m�	������˵�=Uĉ38����Q��+��C����'��8�u�k�5�w`gł�1w>���;�&��yPVo����J��mVX�A�]��-ʴb�%6��^����!�%��n�mӺ�^Rp���9��A���z�2�}͜��q���:��7��F_5	��7�{�~܌���c�#NcT4R;�W�6�\��:�k������tD��n����]�ggx
/��q�ݷÇ�W_2G*-x2��R���v�<=v�!�u�����{=�Ev�{�*C�.�ʉ:��ޟ'�Ò�c7�������˒���{ۃ+�Px��=�OZ�9j�2�J�f]�VZq)��ӣu�+wgYT����dW��tM�v�������A��;a���G���r��8�C�לH�*�鹽���~�zIq���'�Ʊ�W�\�g�|�S�ڐ������Ub���^��
��.c�|l���ۏ_�sT�#`o��뗆%>���ǁ�r���3�Bgh�}'�=�6�.��:n�:h��#܉��;,�5�g^�ݺ�W�N���E�*�k$y<�753�j��;�ű'��}��������|DgG:��y�Y���&�Ǜw<��G ���>Û�oj껄��^��z��g�n�s�9w}@�����v���\������$cn�[�Fo�bA��wݞ��d�ȓ�hFﴦ�Y���JO�On��^��H;^oW��|B@BN�à�>�__�3�+[��}8bO#
����pnί�D���·�{:2e��1�4�r�k��{���x]D�)��<���%x�IK&�#�V1��	TV�Fl�:��^�f�5�X�E:�?p?g;B#	���;~�;|^�yK��'�f�F"`NzD���}�^�5�	޵_tf{�i�C�V�L:r�1��&�L�8�6�P7����S>�>�xXE&i�Dy2.�پ��8ض =��V�r��b�7�1'ªp�Cbu�.�[�+���.�/g!�՝5�@���Ս�*@�g+D��CUPn���.��Y����6n�F��o�[����f�l�S|3\f�;�f���������vws)�P�d��{�;�YTj�F�Vؙ���:#<�p�7�w)�3�|;���X����g��ozH���o���x�ɲMձwBP[�ͅ��u�	-�a��;�5�8Oo�n���K
�p���N/�([x�L*�b�]�r�s����[[��WΘ���'����0�-F.p��w~k�Ww��\Z���Kam��6���� �E�T06��eמ���hM�����o10��u'��yW��׶V&��Js�Bm+<�s��?>+U<�"N>�s���sW놕��'}�<�r���s��Hk����+~�u �z�S7�M�M� z�ܻ��S�{st�I��Byb��+���0�*�[Q�>�����D0�}.Q��oY����]��N�,CȼX��G.���BR��j�|e�����6>��zy�Dl��]��pq����������j+Nr�cB�k-i���ΆgN�"�m]�3l���A8S2u�t;�cM��yie�f�=�K���)�veY�pω������Po��BdÝ��˞��c&�	���>���4u4�&�׆Y�9��;��R8��hټ<�#���Gۙ=��ֳ׼p{_��ܛڛ-dIŽ��)�M]�,ּ߼">��鯷`>�#�e9'y��p����uP&�8����q�(.�g�{���|׽!Y�g&��:�n;����;�-�Lc���:;��>�xi�����U�@7^��5�7��`c�{���?x��3���زݣS�o�9jIL"l����'MzGd�W��w��ת�L��b��<C;��YZZ��;��u��}�c��}� �]������|�� *}�=�,Ag�jc�?J�ż�g�9C�n�[�s[��xΈ��f<�|��Y<�u�k�0g�[Z�c�ޛe���}.�;���wo�|�D��s�6�]+|�Q�qY�gu?lu�<��z{�t�j����C���U��;ʠ�Y�8:3kC��2��pi�&X��x�����`� ��޸����tvhI����W�3^�7e�+;�����sa���k�� �Ǟn�ـ+1=fo��o
�Pf
F
�IV��/Ю�$��2�F��l��7�ު�D��ʬ<�(u�����M����o����}N�zb��ܕ�V@:RpZ��a����×{z.LT��m��Q�`�O �q<�|=��$ޢ��ݹ�6�7�{�T-���<龞K�[�ߎ������S��˃����F�:�y9F�d�5��8Z���P,E)x���kgn���������C�-Aܦ�f���ڣ�#Q�n�jq�k��wR6�!�d�_Y3���_�Źl2����CUޚ"�#s�~Ȅ&�敗�F����E�B�X��h	7���3CJ��q���N����A>���{}�|�����:��F���F�nk���9���:�M�����N�:e��w���o;U٧��q��U��ם>�0o�/U�y{|bcy ��p#/�{=�	^��tS}dԎÙۊgrEB8�-T^BS�,�	�{X�czj�T�1m��׼7�v+q��NtU�GwC��j?hX 78��r��;L�O^	,Nf���]Ԉ�xS��s��Z��^���R��y��yd�9h�%/>�ys[�é����{��I�g�]I�蔼��0���7N�������.�9�K��BK�硹I�J���w`���:-��kg\�ڛ��nL��n?0��ҽ�{(��=��x����	k/r�0.�*�����{�cnZ��9��4p�`���w�m� L^�.��{���(}�{k�-��#�G+���K˃�Z>ɇp{=�8�ν���\ݽ}Tٝ���*z��%��W���<���������Ь�j�J8�D,��7 �;�y�� sƙ�|��{㸛���$z��ٜ�����7����.�*���~�����#�נ�j��bp��wǄ=ݕ�.�Sh0�m�\��)�q
'�s_ F���Z�4iW�7�P��}�/x7���{֭��b��3�'�{�j�U�^|un�jg���D���R�Z��HnH�gd����b/`ʙǳ~GϘ�E!Ļ���瘝�\�"E<���j>��������[4��X**�h]���Q�c->1dW1�l��5�re<p�t+\�\=kq`�6`��p,�]�!�/$���4������Yđ�m]���pjk���Ɇxgp��I����xp�o�uF����)���i�l?g�WI�A�fR��I��rb7y/��&W��h�>m�5aS$q�unD�=ݻ}�=e�ه�_�(ݾ��=��l��9�`�7�?��e#j���l���(5�l��G���{W,�.�19G\�aw)C��Ko���#w�� ��?{7.Op�oq�����`�+�������9�#�%o��'r׻�+�f�-.��Մj�k��C���Y�ʅ��/w{q��Չ˓;�g����/ӇY�u��e��QiW)���ʵ��B ;(����"w<�޻N�C�w��\ؽIVi��V=�qD�����ef�܂�%�\�l�)[o'n4j��M�7�G U5�D�.�u�@.�K�&C��Q����)�Y�ղz;�g,u{s��������l^��\f�Q�+�����;6_]�>6�|��7�z��UM�`����T�o��빫|<��8���E��u�)��y���z����k�nq��.����2���0��c|tAd�7����n6-W^-�ў���t��Ox|<���.���>��9�l�Ò٧*
���ݪ�n�}N�(���4���5R�Η�3�eu!;��=d��ڴ=􁼺2��g=�go��T�d��Kx�o�P0����]ҍ�����ܓ���Ϟ��_/l��
�j'p����.�=���Jt����[۴C����N�t����D��2���7#|z���|f��İi���d�y�\��6�nR�{N5��,x�����t���jB���R*�kXϰg�ZaTVf^��4��[���Y�0�u��B*D��u�:C�[��\#�ꃖ����A�&���n�{=��CWU4.Zob7����:���r�kr$����7��͙�~/t�j�#	O�{�&���w�w��Vo���]�T9�+���vr6����ϥ��+�_E��z����6w�٢v��LtFm��i�*����"�Տ8��u|H��-��onf�Kf�i��}dEv�[�h�_��Sa�����o�?E�~^�����!^+a��������NV;��J�޺�� Y��}t�^/�M�e��+�v{��'s��ut��
�.^� �x��t	.<��N���E&����7j��Hݛ�3l�2���s�+5��5jX�fvǭ��MڼW��=�	xOc)��w�|�Dޔy�^�μ��9t�� �ՙ���t E�I��h0( ffF��f/=���\�)ocl�a�Z�m��ǵl��nS����p�,~��������Y}����_X� u��<y�ܷ�W�L7|wE����f�p�B|���W4��7<D��:�x���A��@�&�����=Ҽ���s�U�;�k�a	�Ҭ-����1[�U���w��#�'���>�Ok��)�����qi��o������쾎�� ^_L����\Ç�2��X@<����)��>�K���+��ΟD��r��gj�O�9<�<W��4*K+T�h"Tš�D@[�̬v�(�>�m��dG�靝^U4���,�
EZ��$�`��O!���2׃>����������Me�=0x{���OU�+Ѽ������e�w Rz�+����|����پ��R�=v:�yD��Fw*kjݻ�����}����ɳ@
�7|�H�01"}�� ���8R*wv�ƍ��H{��Qf�f�e~����w~գ��=WpBnݽ�V��{+E���귙nls�j򋕞b?꧇Q��������P����<W<����~���)��}Fn P�xsF����s4�%����*F4!��K���<�(/��Wrx�hT��a����x,y 2\ҥ~�p�5M����	����n.��f�H`�}�Fv�	��{�݂��<^�3wC���{Đ&
ԕ������+�X�;�iĴE�Wd8�pwv{��7�� �xxmY}�s����Nd�~�e8���ك����y�bL�����j���cyM��ڐ��xfqf��TV�3b�ܵdH��}Z}둥�F65�=ri:�2�S�_x[/�έ�q��̌�3{�n�*^)���:����Xh=�s�;� �-SVؘ��On
�w���&jn"�,��߰3�
�$��^� F�y�,OW?v?u�6{}�\cy��`�:�K�����.�o�[��K�;���ވ`�P;�.�0�������>�f�^R��ܝ|�a�=���&�<Ac%��x�h�N�G��R8b�����wM\Ϗ7�n����M�'_X��M�=�}�;/���uN��h���Ms;�z��Jė_a�^{a�ڤ�=�pf&���O]Wv�bM��^U+�e�<��=�9o�s��(��,K77g;��[6=���*��k�kVj��ŨD(N+�븵��r� +��������������򗽋��|+���{�>�=p9��w�<\�ן� I$�����w���l���q?{.>����k��+��'�
��-�����9@67W^���M�0ᎌ��]�Z���ٻ��n��O�Q���5d}/���9����mq��JuPu��T)�	6���[[���Y�����������ù���;���Gn�#kv�c6��j����0�i7c<�`z�v��u��>�b�Q�4<�y����3>��{I�����^��h�Kl:]�s�G���\�秴�̰��N�On}q
sm=y�ZcslNp�L����@lugb�⃕�c]�;s@�{<p���ͻ-���Ͱ񷶦�w�u��
�ˎ�����7rglX��y�ӥ�ְnn����bC�;�W϶�YT69��Wm�#vG�oNL=qc�!��s�nh�\&��6zy
2�9��v�u$�j�Cۯr������ga�Q�y���ڇ)0]l<����]�
n�%c�����6-�sXKѴu�\�G%^grGg��7���T����w=��u���2��v�/e�`+��<�x��p	�����ab�/f.x����u�l0���-燊��N����5�W7��Qg{M��h�`{ ��6�Y�Ҝl��T��/)<l�u�mg����;8��zj�i5�4�mm��)Ay��a���<�[�"�ۅL%�0��璸��<v�H�K͠�a���G�i�m���uT]�xwQ�\v�u�s�n��v2��ۛ�d��um���/T;��4G��ֺ6���*S-�=�F����=ix\K��e��қ[�����b�>J+��j���c���5t7k5b���v;۱�M��6g d;>]Ιq�(�`�;=)m�9+�a�z��Ѵ���«��������M���6:�޼幖��yR�8�셅v{v�vԽ�����qQ\=��7W�n҃�S�b2�r������X��Y�x^^�I�T��mSnW�����5۴����l���;���v��3�ہ�8<b���=7��t��H�ɇr��#}����a�(�o������P�ri�[q��!��?��G[�&�\��t�=$��|(ǐ��bb�0p��&�����ݥ�cA�c��\�w�Il���fo���a�� O����Y�G��;�@p�(�r�|��P�}\~���W�-�w'B�.7gV��z9��L�jrk>ފ�@H����Z�}���0.��������V2	U��:�����#KNB�9���%�!��Z3�ա�@|�C���81C�G�C{�AW���0����}��2pc��vo��vb���n�v�e�pQ�B�[6���B�zh�֞k�J�}!�"�'t�<C��GI���j:��{�:'M϶��lԱBno����3�m�f��W��7�g*��౳���oh�Vj�8�ĉ��*߉��`�nx�G��"�ğ.����|��צ%4趂7j�H7�r#,�1W_�؉$e�	j!e�
�[F¼V�����e����0���>YK�5�@����æ�{?>�8/�ȎWb�z�C�,�2�c���)m����/PI��`�o�}�g�Ï�(I�%�&�N9k�Ak�+�.���h�鵍<��%�gt��m���(�,��Wi&�"HA���zk>��5�4���0�y�CX���O��f���	üٔ�)�6u�"�r�M(g�c�2�>D�*�|'�"�6��7N�nҍnSq]n^���i�96z��WK�b���{���r��pX��ӷB�݅�'V�-[a.�q�|��v���1c��Ϯ���6�';�]>��Aȷn�۶��;{�Hlt�F�Hd�۱�6���j:ԽZ��b{'ov�gS�r(uϬ�ݷ�z	{7����<d�N�=�nK����m�:��ю�Hk7H�ﷻ{����m�;�t` k��i���{����&G���;xM���(<��x��˜�n8S�x`:4��0��S������"�s����۾;��y��D�J`��	4�4��l+�y/U.&�7��Q�G � ���-n! �p�D�wcW4�&v�+��]�� �Y��wWp���)PnD�ɧ]��g6xf+�����bʥZ>���iFl�i�fa�R*S�g�[O����)��U��j��ӧ7��3�@|��ӄ�ce��.��/��=z�V�nyN������I\�s��f�����`���(4e^�]ݨ��$�*W����ff�j�q�GˈH3�m»�xft�;�u������"��[q+.�8c�g�+�FV�#Z�կ$H���X��Ǔ4�7G]6媜#�������*No�!���'
�C���#�9�a��Ӻ�x6դz9.�e���	ɓ��p�l����i��i�S��n���B�p���ޅ�V���4�[H�-C"��	��v�� &%�5N�mݻq�<�����:zy7gϹj#B�j�h!Ji���Wuo������t�Tx���v�#�Y�}��j$��h���8�XKŖ��wL.�Iѧ۝��C\V���\Jq2[a�a4Ry�l�$�i�S�«Wo���>����m��?�X;�I%��p��&�|7{US���y�9uݻq�:����}�򄰒�M�XI-ݽS�J����Wu;�d��@/9�X1TY�I����1����!����3��<����Pɮ3O����D�n�-0��b� �1ٗ���������K�q!��.NNݮ\�tD9й���Ğt���v��jҕC"e5 �J0�)� Ns��v�y%SMڝ��w}��N��t�xE���E��8)�]ռ/hӦ��<3ckc�*�z��ݾ {��s������⃧s9i(��zݱ���n����7JjlU������#��J���=��)إT��i]��2�t��N����)Qf!�a�Aڻmf�]��]�j�v�y%SMڜ���
�r���P�eF��q�C9�S�U������ϩ~��nȖ���"�>�a�1����{T��u���q��E���tE*�'(��E_OUd^�A;���%��w��N�Im�T����U�ͬȾh`�Kr���qn�n��N��h�����Ho����gVO7;����'���)�����@4h�(��$4���'y��B
�`�YA�eS4�Z*�S��^iVn�j�v�fu%SM�����(PQ&s����l�vۇ
ݺ�}wg�R��s��½cz9Z&�K��Fk�����_����osJ��k�<>�\�ήJ��R5�r"T28O��ۻڪ�Y�g[yt�)���qֈ�|��:����BA�mC��e]յ��t�-K��Ni�ȿ~����@���KIH��jU5��&q���T�N��T��iWu}��K�zͺoR<P�P�%�e��]��j�S�ܷ�2q�L�J���9�S�Y
3&gVH��Ff��Y�7��E��T��0.����-�n��p�~<�w���e�n2�j%�ט+$�tnb���(Os`��[��Mh���/z�|�ie��ql%NM��&�e�s��;9�����Dx!㗧l]hݭ�
�3��GF8�N2�,�Zr��V�+��[���y.-��[ ۰/X{[��0�0�dq�'[Dg�:���nz�s�6�F'��m�żxglvxƦ�[����_u�o�ۥtsa��kӞٛnڸc<��Y�v���N�u�k�8�ێ����7et{*������k�z���^{'߳2aM�]�f�w!	���8�������ͳ'��`�چf탛����~;l���v���L��W���W�F�ڒ��=�
q���U�[X�ѧM��^�n�Z�*�,}�D6�m1A8);�Q�I��s8�`R�x�DR�o�L��#�N�Z�܈�&c	�L��ј�${����>q��;ٙ6㧉��m��hI2J��0�.����S�)R]�y��îaO}���{��P�E�D2�jh�ZRe_fػ�� ON�����)���| շ��H"!
H�XH��3��n{n��[ddRr����x��{]N��u��IF"B)wo/��]��Z��A����N�����(T���"\@FE�i�S�E��iR�������tX���$��UM��{Pʸ���y�ې��X���e2D2y[��1z��NOs�������ѰZr��{9�7w ��)�Lh�J;�M��h�D�IMA$��d��Sw^�/�v���Ͼ��"�x�&2
0�ª��X���/ffV:~&����v��'J*C� 0�Jk��NV�ݵx�pE=��]����� �4�f�0R	�.F{91���M7`}��:1�=S�)U;��Wj����IQ�( Y�{=�iy.ծ��x�k����j!a
�8��PbHm�ݿ7����ߚ�]�[T���}�k�s�L�${��"m p$�f����:*��}�;uoOM�M�͋���+2N��ÂBZV���(��D����=��>%�,z��H��@��{�N����>�c��:�?S�|'��y��}G�k�{�DS���<-�f��~���1��sDl�A�T5f�gF�����l�w�I�]����K	\� D���뾣«W�~�6D+>%�n,EhCJH[/�����Q#��-v�z0qfv�_Ϻ7fH�g�
���1��F8���5�O�f��hW�:��y�t������rd��;�Dh�M�RN��nަ�7$�t��粢��v�.+��<��
\AM��4�P�su1J���n��px|��➎�woOT�a�Sl��,�.�^V��| �����)�g7�v�g�<':l��}�`�M�I6cm�v������;�����z��;���_��-Ȋ%0d"��ڪ�{����UJ�mR��C.Ӣ��cJ���]��𛸱�pcu�����ٔ�
�f�qlI���#�����M,�aq�[:�v�c��j4�b�g}y��}_�L���"��	&H��L�LwrMD���o����n�rF�58�^N�U.t ��76�.\#�nd�tn���V+�{�	�!�a1�	B\��6�P޶��8�!ٵn�^'mF�m��KGQҾ%o˽����>�J��lw�}��:��R�{�"��a(p�j)ѻ�k�]��M̝�}�U�x��� ��$��f���M�SM➎�wo�U�s���U���ɒs��I$�(����I��w�U}�.���U�v��ڦMMw�	�u�ю���'�2�0�"	���^V�wV� �W�*�SőTj��+;xm��؝���^>r�;~��h�" ̕�ٱY��LLl��u}�/67	� ΅�3]N0�uwt\�&��i+u�&gH�mn-�w9t�-�X,�d�P��;ԧ�?����o�ͨ���X���Q��%��8����؄չ����0��n���c7�zK��a�4�s`��v����i��'c��ԑ�n9��f��\�u��vm�������腸�\磂NЦ�vwO��y}�oc�m�`ۭ�:�#�$8{�ܜ�p�a�R�r0n�m��%\n����\�Ӷ�S�5���l?=�;�ca
�H�iJВ����}8�n0�lN�@�ANn�w�����w]��>�ķc�e���f��ukK����~���&�J���U�������X�O�m�B�+���i�(�RqN�9�� ��37�v*��ڤMw�W2sl�M�)��)\[�z��R�qyZ��p���źl�
�Tɹ�&`��Tf�ﾜ�}��uR&���zv-���};3��܇�z���F��͏��t�}��x]��sMQ�wʶ.ݾ���?~�d'n�jF(-���{�7�,����n���݈�m�h&����RL�B�RD��y/�E���tE*�9�w����Z�TS��u#���)�T&�l+wm�ҫ.�m1fb�+�5ۛJ�=.�d,^��t�~1�y��'�mǏ�=��gC���f2�����G�6��eWR�43pV֜P���ɞ� D@�~)wW"�(� R,��;]�3�Z�S�g8���j���gh7o�����Q3�D��4㷍�յ�UE> }s'x]���iTs$���[����1��ݛ�*�{�ҹ��_r��)���|$���ʷ�Ԅ�A��N8L�o>��;Us�*���]b�ۍڤMM7�����A�����"v���q�p�.cn�n���엊[^��V�e3D��i���ǫ�"�S�y�]յ�U���No��|��"e	d���t�Vػ�ӓ�h��o%�!n��ڈ��w;ðL�6���i�Wumj�B)�f�E���𜮭S�l�A�j�ؼ�)l�V�ӈV��z-`g{K�;|��_b��	��^�	��{�3}�!��ً=���xK� ��$<f��N��oL�S�ķW�˔���>����rv2
��L�͛�e��Z��w������s�kʳ�)�7�Qf�m=#����D|��G{��ů�8�]\��ߚ�*��d�K����c���7x�f1�q��f;��N��F�'�]ɤ3+d���K���8%TD��G*�{�T�=����tP��B��@j&9@[rs`�U5SCX�2�Gp	�����Ԭ�;8����+��8�bZ����V��̉�9�Y}�gpW@��R��/:���Q�]�4�+�.Ďy/qaSǋ��S6�y�N� .�D�������3ć�������O������I��D��q�n#��w�Ǫ��ʫmB!Gt��ڈ��k\L�n�,w��xf�,`��֘��������N�$5N�o�_Ѿ�&�m��^6��e�ۺb7s�-X�pw[��{8�g읗Ƕ�5%`��;��ر�۽ĥ[^;P��2<��L�^�,��[��ވ��S|�<[�J�8ܬi&tYn�P3B�<¿�b�C�:����yFE��L���ӣ/Y��'�����^e9�F?y̽¥��ʐ^r�=�i�,���sO6vb�](�V&\��r���X�!R��&���!��S�gj���(T7��5	3���W�aѭ�Fs��;�eEQ��x��ؚ���(ӥ3�;T����=�!�s:�p��vb�X�sn�5[�~qN�� )������ݞ6`������M���2���ht�"�5�p���>c	(���#�i;���z��g?k��@�*�wN��5X�4&i�Ð*��I�4x�����Eh�>��}�>�{��.M�F�~z��$#6���8n��V��s��2>% 2��ot4�]�v�"���ԣ�u�P�c,��M �#��;n�#����>�Ft3�I�=*�7�;@��aa�b��u����t�������ŀ�0� ��]��SE^��������z���!��c,�־�$��$��
9�N�"��I{��ı�s��G%MӸ��m3�e��*Tי��?k�,d!���8b{�5�Ӯ5��+�gp1��0n��YLk����j��9ԏf�^�q�^\1x��tfv�y����k��F�3x=�p�T�����؁o!!��V��%Tc�6<!ޒwg ���U+�x�퇵q��yw�\��`�"E��ub�6yc]�m�cH�v�-�Ա�h�+�i�㐌v�$��K`�j��0h�i]�!�貉�Ñl��1�'��J*Į���	���z��[���l�|5jAkޒW��A�} � ��c�㋃�^�;n`@ݚ�i���<�s�tf��}0Ѐq�(���BR�L����y����B��2+t�&.4/d帴���`��J�g{2�p��뤆�
$݄�bB�9��.�s� LT��"�p�(�h��u�
�����.���,�~2�Mr���������^��q\
#���M�ұ�e4� ����5�{�%�{��v���L�|i��_9�7��3i��+��hj�	�s�$�~Q�b]q���L���'���-�H��9υ���=�cJ��BD9|�X���!z���_�Z[���m@�M�Xh�)��{tA�{k��9�͍�z��Е1ŭ�[����_m��փ� nt����﮹�4���26e�«��M��A�Hq�9�l�M�
гP�߾ ��BCm�8��il��ֱ��i�Da i6��㚿{ͥ�{��v��L�|i��_9��x
t �}���E�"�Q��M&�6i��e��9����7��gk��g�IUP�VG��n�a�y�cJ��BD;��5I)�FKq��4%UR5��(=CB{��u�!��E��E�
ƚ�4���x�m.�1f{�u�s4�$����ě���d&֪[�z&�w)��rw]=�.�g�Q�pl��.ޡ�#�,f��槺{+K��rW�l7�������#&�w �`M �/�j���~��k�B�7�FPD���ӳL�~4�M�����ųim��w���l��)9���.i-�Jf,�a�GhW�:=9!�f#"H���I5�)�n��i�(���;�'��֖��{��:��$�2ԍ��j��k�,��^Ь�-4˿�s�7si�o���G��$��C����=ˮq5�,վ��H�q��(��+k�Whrgz��� �2Ϲ�gk^6��ƙi��s{��\6j}t+k¨��#���ߛ^	8
	��.8c�a�q5�^����L��k����Zza',�����0�5v��=�.�E���_N�(����0�cq0li��i�P�UCy�O���!��E�����qV�Y�?��ˮ��ώB$�Y�gtm��ƙi}��q��QJ�l�ۺ���G/��ڱ���5v�$$�����Ķs���|4i���2�g69Oل\}�&>u'h��D��&z߄��G��;QK+)�!5�4�����x��FD�<�Z�t�j���O�����̍��۽�,��M�8o6~���S�N��j�$��;:��a��k��h�j趪�y<V�M�.o������=��}�}��%���6)�7s�n޶鞮�(���u]�p7.]���]�d�+���vx�I^��p��;�6�p�/]��rNE&�1ru�m�6��t�����om��������,n�S)<��r�6�[�0Lc6wm�i��������ڎu�ٮ_I�c<�9�)�h�ȟս�r���x�ADQ�r��2�ЃD�$D�7v���\mD,F�O2�U���E�۴7�λm.<{m�[#�s]��{�VK�1��0�@�j@�~Y5v����\#s�Y����������};�? �'9�q2ϻ�k��3)�]�s;�&�!��Q��nn�E���_Vz4i��{��2�g�}���ƙ��Wk�h��2�L�����w6��d$�>�5�b��Q5		D��X�O�V��k����ٴ�}��X��i�}�l�~9Z��Kf��v��IZռ�ݔT`��lǻ�窀Ta��p+6�M%�9�Ѵ�7��g{f��1��>$d�����s�ٴ�{ƯS�V>��R	��q�cMaj�L���p�5�"�@;� 7�eo�l����ع��h��S軡X�VF��C�t�x���x��<t��j�c�ex��Ύ�J��+�m�xLO�t��{�ݾ���6���*�,�>-����Lƾ4�Nr�����l�[>�{�c�<A�M�I�g?���s�Y�q|p���|�[4��M��E�� ������T���̍��bG��� =<��G`W-�aÖ�]9.1���R��+4�Qn#������ч1C����(��T����_;�b��b"�����=t�h�-�m_
�3^ȷB����5v�����k�B��l�g��}!/�f��{���8��J8���,��K��nƚ�4�#���������Kg1�-e0�f��S��CHf��"�}��p��I8,u��|H����|n����S=�3Fq�]2Ӝ���Jf�d [9���l�4�!}g��D�JI!Q�ن�H�ZE3x�J2�L��I$���6�fҙ����f�i�R}�t��&Y��zK�|m�0Tq��fղ��1�=�m%:��"�,�u�v��	��A�����������t���p�#���_�֑i�/�3I�Roǭ��m2ͥ���H0�#Bs�� L�#l(ڑ;�L�IL�+��O� L��i�{�w4�f���њ2�&YI���擤�(
��E�W���*F���\0��v4̦�I�__74��%3x�J2�k�w��:z��gʡFֲ�(0��>�zr�D�őY�6D-�t:�{)I��O~�QZE�Df-;�kAΗ������j���/���(���D� R(떍p��ƃ�u�x�!=���0֑s転ƚ�4�"ru��S���Q2��1.��5�D� (Y�v����j���WZ^�_�o3F�Č�NVz���٦��������L�ر��5
����5�C�D ���m��e'��\�e�J5ߠ�0�#B< �u�0��	��t�r�'<i���`P�����e���6��	k�0U ��n���MG#��3\"�/��,�2�e&�|z��[4���(�# e��i�o��4�M4�_}�8q�h��Ԃƚ�4�!}�F�i�"@4ͥ���1FS�s=��4�f�\��ݍ5� ��pՑ�{�	�HH�b2���"�i��� �P�5U���\-:��������f�i�R}��m֑���k��a�B�`��J8���� �=�ˌ4�_y*�V��u�W4n}�����wP��Y���7���/ұA�>Y�Of�ٞXQ�^����k8@�T^١&cV�썹���jUk}�[�e�Y�P�Ȩ� (��x ou��qxuӸ!Q�J�"-��^v{軣f=�����̜K�*�e
T���pF�Y����'.�v�5G�mu��D�z_nwQ���+mWi����W��[�Z�եM,�Z׼�:Vvb%J�W�����sk���B�.��0L���0�(:�Ku�> ��r�{ݨ��J�����tP�UC9}��|�W�q�/{ʦ��2%���� >����I{�)2�&�x\,j[�/;T@��-���|��~^?Lz��m߅
�*��>=�7i��H�_�)E-4�PX�VF�����W4�f��Iē�H�{F7s	�Rs��SI�i)�n��b�3)�Rk���F�b����c�͠�[+=79�,���d��=#Ca������=�)&<��A�R�R��#*�.�vrh����+�b�;�M�P#kfq;2�B`BL��6�Nq�j�q��6�B9��yۻl��s��\>j�[�Wg�nh� [��ݹ@\�����f�x�sE5��燵��l�k�C����;/R�շ��K�e�N^�V8 �da���j��-דn��ӻz}����nvx��e�cm���kc��\�ۮ�Sn-�k���mv��	�s�k;�x��Ϋ��V�1]��W�g��;\�=��{f.:�$m��~�q�bۘ�dF�h�,AF������ܫ��~>����K��Gv��ݺɷ��ۉ��x��z�U���{��o�펎�ۛi
��w{���w�|Gg�TTe����,�����Lj��x~��&Y��~X��(��HHfSL����ۭ#i���G�@���Ie61f���)7�������6ͥ������>���&>.�7��Q @Yj�\�ރ�2\��cJ5�F{�%e�YI���W4�gH�$�&��~���L�e���z��i�Jgտ�T�Gh�a�Hݍ5�i�hUT-9Y����٤�s�іRe��V�~wZFoj��
~�Z6[>��p$��Ȕr6f_�H���a���jUQ$!�k�M�ٴ�}�ﱋ4̦�I�_OM֑f��k��U��n&Td�ŉ�\��[�w-��Z�[az;�����{k����x -HnH9`���c��5	�s��sI�i)��~�FYi�R}�q՞�0��i�Ke{�b��	�RW;}\:pHE���ikH��/�7cL���`~�7����Df��UZp�佞�������j���3���C���*�K�:�
��^������M��2Nj�{:��rM#_u��&�F�T#h�Tlj4��qQm�k�sr�5I[s�}�k�Ʉ�g��Kf���w+FYI�R}Z���< �
�\"�}���a�RKF+�i��e'���\�e�Jew�b����4�M�]jm4�%3�_}�X�XF��r���n�3����Rٯ |Ig+�Z4�L������,�S=������/�!x�z�w�H���!��HJ'ƚdi�G9��4�f�����+��cm2�e'1~|��[4���Z2�L����~����(�c5;GŷV@�vyv�oj�vc��u��n�v��7?��z~���Ĉm��F�ן�0Ց��\㫚L�IL�h��H�I�Zo��+H�ZD5މ� ���BCq��3)�Ro׭�>�HY��s�іRe��V��4�f���w8h�<@��VG>ޢ�Mb���(ě2�,�S=�3FY��)5���{��X���rJr��P�T�,=�K�mDL�_VQ�<Ko�k��O�=Ds}p�B�iU���G)�᱐�,��8���;;��s��gZ���9�'��6�
I+gv���-TZ�TQ��F��f�+r�i��o��~�,�2�e&�|z��[4��p���Z���(�M�e&�@%�/�}��L�IL�=�4e��e'��\�e�m>�B��Y�4�&YI�o�#ߜ,e@ː�ikH��/�7cMa�@1$!�ϟ;���_�2�L������H�ZD5�U��"���$Y�2���o9��MغP�+�.�k2���k�Hۚ=r�_�{ޠ�"�vmG-4�R�Y5_{ήi2�%3��4e�L��[�<I$�M�il���ci�M2������X�Hʌ��7Z|p��_<�� � Zi��^��4�f���{8h�-2�O�����#$��6��c=|�XP�!-4�4��P���2��5�F}��~�L��"HCl��3��ͥ�Iy߁�B0�!o��8�h�j6���H�[�� *�zg��MYjϺj�,�S�ќل�Y�bV�o?Q���y�"0*��L�C7Uo-�+�E"è�[��N堹���ج��r��\�,��M��B��y�!�d(&�$k��3ma�ox�Jb���d )[�nF�F�U�F�sU͹]4Rb,c�|*���ύ����E�S�Kȩ�5��i����4̦���+>|��[4�� �@�o��i��e'վ=��&Y�C^w֠�VF�xUߺ��TbN�;����b�6�m�۞x8�;j��x��d��  wl��
���f9��,�S=�3FY��)>����,�S>���Y�f�l��/ϛ�Kf�y��1�����0�V4�#MB�Ǯ�O�  i�g�<�Lg�tf^?�݃ �J�
����I���F$7ZF�!����ƚ�4�#�:�ni-=$I	6��f�}F�I�R}[��u�a�"���1��M% ,��X�Zi� �	-1���ͦY��{�f��	�R}���&Y��$> ��|�p���|;T��`����Xi0��t����a�"HLs|{si�p��j5f�#���n���X�r��������gJ-�{���l��h:
p�����N]us�h�zi�s;VEd�/��y�$�3�`��l��X���M3�K���?~����߄�ْ����D�gs�tc��N~���w�9�NA�z\�;���3|&�r�,��H��"��T�JRx�<����V�G��M�Yy�։����p����j.)�o\�1q#����[�Tb�V�AV�x)��vn�7W���L�G"�Cqmh}�Sy'ND=��@��S������76O��'X�括�$��5�GoVD:nb�J�^�k�\�_��R.tPS�T��&�'0Sޝ�\E	"KW�D-:�)�޻�i�����!
��(�F%.5UM^� O�"v�p�E˷}������E���Lu�~��'�O������<w�����6����o��^��m��+�x�:簹*Gu�6����;/���az�YG�tv3"��"V-�$f���uL���=�����p���h�� 'C��+�M�����r�?��2��K�/K"�r҈3�e�T��蕰�D6�m��Z���J�*�L�v�t�d����wQ�b�jG\��J��Y?u�Z�u*�3��� �=�y��!� 5�n�����Nާ�˷�y���7u(J��y�g���^@���{*�2�\m���Qf�$]�+&TY� �uxb���d���|���x�����fY�#�Q/3�K�yN�l�nj4+�w|�����7�\,�a�ˁ�H�&hmt�Uj����n=�{��ћQ�x�݌�G�n��z���GGOk��<7m���ݹklc��]q��c��vj熍F÷��@���8ƻ�����;�n6�x�w�^���8"p�X�>��b�����Rѹ��݀��F2�"�))���&�m3�;�3)Z���f���뇫%�^ۻR����$�����s������7�5�WQ^:�;��ۈ���[=lvgA���:6�]`7%�b4-5�)��v�5��v9����G`�	���Wg��ˇ���w7n�	��sh�������vݶ��'2i-���t\�-Ҁ���{nt�p7-���j�$�<^�\�u�ms֦͟s�c�Z�v���#G�����Wv��o7}�� 㛧N7Z�בG�Ϸ�qTk^�7nѽ�|싐Bg�\�Mm�Ý���c�]��A��wFNcprWlcW1c7j�����.�<=����h�b�Φ�7�{c��;ݹ{���}�]s��0Q���s�&#qú۵�¦d:+��=�q+�ۮ9,��h�V��,0�
��ˑ���ɍ�(.�t�oX۝��.7����C��m`���n��Wp���3'.=��HH��-B��;[I��'<��M��N�2�wimv'(nj���Ue�����:�R*��c�lm�g-�����Kz	B9�^b��Ǐm��.�әj
�Ng�q���0'<ڱ�k8'=�ʭoK�:�u�]��ݰnf3�$\vS��JX���;�D��2���y�[v�ݶ���Cd�g��S{�k�ۃv،f՞������x�s�c���M����0��3du�P9g�-�ݫ�zv� h�z�#mɶ�N��;�}z���:=i�����՞���0�g��W[���n�d+B�=��{r�:Lݻs�z��ͻ^�h8'�v��Kd�(;��NQ�󳗠���ㇶnͣ����l,v��̓�s=�:������٪x��-�nۗ��9v�9�3�k;]�l1������c�k{{v�-"�w.�e�:眧��6���[�B#���n�}:[���P," Ä+��1#����L�S4��2�æ���s#�F5>s�4�85�P�مf�0�#���͍@��VH[�-9Y3��az42�;��ǐA���Ȅ���=]�k�[��>�h_8�!|�An��!�|Y��Z�(A �`����՜"�`v�#���|B�4Y������E{���������4N``�	{�� {����w��'/��G5�#��B3�:G����� �cv��\B�z�ܰ�H���Q�|V�6�+ڇ�ٻ�:5��[������~r��2Ú��#���Kt�0��p�S='�>8O�幸f��y+�eDO��8@dۧ�t�>�^ d{۞����� T����!��;��#���L��� w��nk���<Q}j�F��W�0�*��0S����L��o�I�>�r�p���&O1O�S	�qd��os%�i�x������i�����h[���c�k��;Nd��ϕ���B�_4,�D2.��C'sQ��g�0ǁTh n/v<���y�1���$C���'Z�1��3Y��o)���8�$uV�V~hHC-K��lt^on�8����6c�s�yصF��I�7����X�ɺA /JS�(��?a�'��O������T|�'�kN��
&o�_& ��O�9D��g� |J�&5f^ѕ+v�[(+�/
i�H�q�H���ߟ���rlQ�Gg�t�7ަ6G�[�N���-+�3�f*�g���Go]�d�Z��L�������9�2=mp�BZ@�[Gk��y�������D��7�����v�7F|�ۓ�S�+{`Z���[���y�D�x��%�Ճ��{y���pL�`J1��BMM8�&I#p�]ڻ����%˞�:y^s�auZL�W����qˤ'���n�g�{��������h1QXԛX��kQ�lZ#%�X*+F�4i�j�ш(�nlmE��RV,Z1�w�z�����^�yܜC�n��9�9\lN0`5aK���+�y������J����Ёbq�R���Dt�O��{W�L�;��fXa�o�u��$d���!�I�E�d.t}�
��D��j�,�}]��[�FBaI���i�������l�}�s�4� i���:H��Q�ؐ��n��&����0�a����C�Be�B���p�5����PY�#�P��|�E<�2c �L]ik{T4��
�z��L�u��w��sI�i)�n��b�3)��AKNf����Kf��ޙ|��_W�E�4�M2����i2�3�	'�Y�}f�l0��|j�,�S;�24��P�
���j"
jT�4Z��Xו뎑�Γ'qCum�v	����uۮu?�{���[,���p�5�!����٦e4�M�s�4��%3x���2He�����W4�I�}�g����X��mI���4�!s���~��C���*�'�4U�w���t�D�y7?@y�R���۸�;���7,�ȋy�}��t6�i�3���kL��.�@?|f�9�����@c���F�d(��\�$l�"�d���1QƢ1V1�#Q�QcQF�Ab"6���"`�A�1hԒX��(z�ϒ�����߯�&�,����+�B�4!�g��#�2�n+�0�a��xjKf���KN�`@�s�}f�i�R}��W4�f�㿺�n�
�%�����|�%�;�y���4�Ϲ}�1f���)+�
�KfS�	Kf�=4�L����*8�h�j3�ZF�!�}]�6i��e>$H@1��w6�fҙ�Q�2�&YI���74�I�t&=}�ғ/�Jă�[�l�	qՐ��MS����`I�`�7P\1��_���wG�|b�u�tC���di�G�|Ĭ"�aֻ�1��e'���Y�i�m-��{Tli�#MB'g���J�B�fI�ZL�IL�h�}$�!I�Z}�k��&Y��}�ﱋ4̦�IX�qS)貁���ij�:�a*����1�����j�z<5�B8�Ν�)A�us����ShG�k�.¡T�>����E�����ᝪ_t�WTa�X�
_DT��Qq��_Fefu�dt�zr&o[��g�,�o﷾ίwz�I
��[5�%�5�Q%�W.m��Q������6H�E���TkQ�Q����XI��F0R*0<?9�y��7�� �L�!���p8Jh��r�M��22HS�_}�]�Y��;�JfXk���l��`����������,�N��n4M�F'0՚0��3S,2�zH�@����a4�O����,�S>���ŚfSL����{���ܵf5���8+g!m�1Ż]�7Ps���u�[����j��w����t?w�gr��Q_-V1sil�S9��іRe��V�s4�f���s�,�A� �2�e���ۭ#i׃�!�L1)DPU�fa5�wW4��Hm)�r��b�i�a>�}S)l�}\-��	$��Ր���!R@[�Bl�u�a�%3��Y�Zi��o���&S�I6��z�Q�a2�O����,�S9���D�J�4#-��5�i�UU@!�}�M%�)L�/�FYI�R}Z��L���.Qg�ߧ�Me(�}w�K.O�[�����W6����v\���"͓1�h��OLR	�?]*�9�;u�A��)Ќ[�۵�O+��n�ΉτG�""#�lb���&5,Q��EQQ�7�F6��6V2AQhDB,�C�$Y���Y�Zi�G�ΤJc$D�AQ$ĺ�,֑w�f��	�S��&9�u���6�Ϲ}��i�M2�x�w�Kf����Y}�9��ˋ�Z��C���mI�nj��\�61��.I��~;��_u��>��ѭ�k�6�M����_�e-�Jf��h�L��)>��Љ i2�%���4e�L���%K� c%-Hn��5�C\���Y��	$)6�O���.i2�%3ؿ�{¯����m�|Aވ��-��ph�VF��/�2VddU>����>� ��7oѓK_zU\pO��B7Q��WZE��U*��k�<�B6ϟ�)l�Rk��gI�:�Є��ٚ�5e���ۀ�K8�e60i�F��>���T|x� �;�,åw����J��Wv����4h�Q���[Ho�igUa83'F�N��*'t]W���UHeTCŢ�+fv����U�кq>��U��o��q�l1����d�9Q�uO���s� ���w�^����B�ٽ��y$���ֶF�O/cU���B�V�uC[4BFF�M�z�+�g�Z5���K����Eܹ�=����.�}�`����=�m٧�n������i�@m��zD��j��Ȃ�l
[=���+;"�G����mA���'#q�;c�tAvV�&�+��0��[8�v�a[��$s5�0�����n۷wnX�A�����͊�60%&�+��ђ�1Di�?��r��]��on�lه.P���\�4�g��/!p`[�����}�ܱ&MV����=��Fh�r�c��x|>�[�ӳ�H����RHą6b���ŏT��<P Vr�Y�m�/���z���� Vr����*1!e�#(<�߽�ܛǟ{@C@t�@*��o|�|������Y�"��g��
A��p�`��Q4���L_:�6�f���w�5Y�)>�L��[a$!L���(���w��@�*9$7A���s�c6i�&��� }^��2���o�i�����5�3]�,y���rI]^��m���Խ�X��.������g.�*B������{�O��Y8��+�V*Ͳ�l������9�e�Y������ B���}9���l�4��w��,��PCE���f�D5�|!��wPg#���WJ���R��zĺiՑt�U�����>ˮ3��k�9�z�a��Y9y]�{V�P0�����]���i��VkaQ�(��W�h�X��H*���HC��)>�i��R�5����̦�i�:f�SD� �i-�gˬ�\ ш5ƚdi�Gݙ�sIL�S7|�3Vi�}$d�e���r��5�C\w�`�P�5\��a
Er(Ai�u�Y���U��~�6�M2��t�L���1�l�a��Ro��73)�w��}*����|W�%Ӹ�z��5�C�@T93����e'��T�[2��c}�f�i�Rv�p��.(#,��!d%Q�:Çk��V����nw\cF�d��MqV��w����닑�I�u�,����a���j��x��S4���=�՞�@�e&�iO�r��5�C_|0���Da09��Ri��s�je�!2�%�x�vY�Zi��s�je-�Jes�b���B4Ր���	쑲�@�K*Cu�CZD4����k�A��ī"����s�����7�J�a��x�m8-����b�}"�V^��ΠE>�\u��8��r�����	����}����;3�]���AH�DR)�D��AIdGЅ��|2�&��+H�XD4��}
d#$P���آ�2�OH$��9�U4�̥2��1FY��)7�ϛ�Jf��|�,�lg|ݎ�4���,G$e$Rg+M���o2�,�ЂI�p�M%�IL�9�i��e'�ᚙKfR����m�%�SF�ǀ����;^�(]��Ufy�=��l����e��㻻�_����u��0bͳ	�Rw��74��%3��;�Y�e4�J�>�G�&�,�[7��іQjϽ��Q��R�Q	u�Y�"�s�,��e	�'ɶZ}Κ���e)��ي2�&YI��|��vH�[6�i_�^e)$bB�1C��k�P�����KfR��_����M2����M%�)L�9�i��e%n���8���!��֑f��B���W�`pk0�e'9��4�N���ﱍ�e4���E�������4&/|2�{���ra��K�8p��\Prč�ɬ���px�%>�V�ɪ�)o����w��S��W1����s�w��>��V"D`�a�1�\36�3�������2���w)~���88�64��B��J�ㆴ������{e��I�:f�Rٔ�T�,pa�F�v��O{!m$ȍ8�h���*k[���lj8M��XЮs�3ڊ���ߎ�~2X1т(�*Hٺ�k�CK���i��W�2�̥3X��2Ѧ��9�R��5�CS�un4
n7pV1X��2�L��|3S/HL�Il���e�L����k�M�ٴ�}�ﱋk5CH�#���@Y����TṤ�i)���h�)2�J�߱2�N�	Il�9�m��e'�隙Kf|�/�2(�L�hG���zH�Zw��Si�i)�r��b�3)�R}\z��[2��@�n�ѣL��R/��;����;�#i�g�e��O�9�U4��%2���Q�20�!s��u�a�"Ϭ{<8�"?w�����Uu&t�E�Wۻ".�$�5�9��3�s���NL
���ێ��H��ܳ{�v����584�t�ĭ�#���rb��󏞃6��N���w$��r�<���5���˭�р�ƞ.`e��c���s���m����5�sӷQۃ�7�nFٱ����'Uuٳ���F���5�5��X,0�S�e�m��7}���ƺ�{Sϗg���Ύ���bq�H�����T,' �`�v5�1\l�Վ�7lc�c�Ů��{Q���4�[n����n(�M�m�|U�
vMȚ ��� �TA �i%�c4�M�лi�����S�3AӺ��3���]��+�ۮ.n��s��y�*���궷ޭ�F�B2�q�5�i�B�>2��5�S5��іRe����>��D&�l�[_;5di�G��1��A�Rb\�[4��;�1F_I
M2��s]ni2�%3�_}�Y�e4�O��Z�O�f���{��d��a�����L��)+��ح:f���_;��e��$�->�MT�[2��;�1FY��)>��))�
)��7ZF��R�Y��w�śfSL�������e)���h�)2�� B��θ���4�Ͻ�s�t�qB�H��5di�B��%ak	O�$���LQ�a4�O������4�ir��v4����=;�KM"K�r�j�:۞��e��+={X9s�+���W[`v�RH�T	a�l�K�I$���6��b�4e��e%s|qSI�i)����Y�F ٔ�->�L��[2�ϫa)��P@Y	��i�F��/��D�q��זnߥj*���qF����'n���u��7e��E`��m^F�47s�=��:&
LX�7�"]Y�柪|#��vo.g��.	h�	 �$f�1�&�2d��
< Kg��׭�i�M2������[2��b�4e� HHZi�G=��BڊF���֑f��k�}��i��e'�隙KO@ �[,�l84�#B�{E֑���j>y�����
l�RF�i�#O�Q� Y:�ji-�Jf�ܭe&YI^��&S,�vH�-����Y�Zi����P��0I����H�ZD5{a���j��+��˚L�iL���ci�M2�?�L�"�aרW��#)A#5q�Leu��V�7�}}�vL����P�7[En����Ě�b��M��a������������2�fR��^���e��I��h�@i2�%����Q�a2�J���k��������0֑._�nƟ 4�e�3]�͚m�Jg1�e&R�\~��t
�i�"�_>�ڈ$�n0X���5di�B�|6�H�ZD5{a���L|�fuq6_���ȃy1Rv�8��/r�T��o��zt{ӽ�f�]H�52�}j�lsSmd򻎅
��]QJs`��-e�)eX9J����/�C��wRn<1��z��ε�y���V�������v��vNߑ�S�ծ`J���۞���'��`��U��^��Kw�l~plf��}.Zx�k���!x9,�]���3��P?[�� �:�<U�}С��l�[���P��:��(E��-�q� ��(���L��L��r�frb��kݱ�jn��~`R�������:��^�{|�^�],��0y�A�IM	~��5����xo|�o�}�A5~���#v�7A),e�B����2ƛ�)6iLlNK��#e����%�,���G�%1,�=0eͼ5�5X�WU��>cg/1&3��������=]��W2��є�D�z^+�9uaVM�t9��{�� ��$W}m	��C�i�ya�o�o��q�1���Y��Иh�8Au۝�f�{_�o=T�M�ۖ6����$�xxwr��H8S)��5+�Tn~���7�L0�4<��U#)�ñ�q��)�"*H���n��l�1��l����̮�ib�J�K�k����A�V��L�wxA��}�<��U�XZ�A^l�7F.����{�~˞�s�N��ѕ�Xr���*V�L�9�Z�؍�˚���*j�]���g���}��2]�Uݜ��F' 4���Gz)}������]q�7g�䜧��܍����ݫi�9xF���2L
��L������7hR��j�!%?(��3|�7���F'vw�����P<3�{��9�PLu�o��,�%ã��55��Dg������h.l��d�~���8^�#9��ZA����`���A�/�doK����۵ah���3��#��xa��;�@Zxzd���˞��/U�H��dl8�kM�[�.!�����o��,:�\���6¬�'dƕ)8�j) Q���P����ZP�"TΟ��X����4�j�T�-Mf�&���D���;�׽zvG3�&�f���y$#� P��I�/,#��s]&�c1C�޾�~X;ۡv5�f�yƳdƷ;"�%#3@�'xl�����Q��7H��j("C�x��x�d�ë:�V!K	���C�8K�|�9���*-����p<҇#�aW<���	����C~�N���"�i�uH�xn�3rh��q���تnh����}�pL�[8S0v�(�_3w��W��g
��0�&�j�\V����p����Q��d�%⚘���bJY@���%H��i�*�H>�\Q���֘�;���Wwg�[�³����\��u���ҥx�X�kӿr�l#�|�9�x�]>�V���Ч�K�3K8� �G�f� �I����	)&q[5�/G3��͐�CÍ�2��̆i�s�١�kHSX���=}��O7�5�(��;` R~b!b�f`1UTE���O��蹤�4�Ϸ}�v4������#��	I�֒ٯ@�&e��mh�)2�J��L���k�}f�i��A	i����l�5�C_xA�y��nEQ"a��XM2��s�.i2�%>�c�ﱋ6̦�I˧����i����a��|��;��r9y�K99�Y i�F�'o]�u�#Rf��{��1r�|�sh��v��!��7)F)�\�a�Jg1���O�)�Z}����&Y��Q�Y�; d�)4�O����0֑w�&�Ԅ@����m��i�M2�wO;��> fY��s�іRe������L3-kϜ����);ΐ|�
p��E1u�Y�4��pY�0�s{拚C��S>�����e�M���CXh}������q(K�cRq�����qSI�e)��3��2�L����L�I����=����9��z�/跋�t�US,a޾�����]��t"��gP²�j���k峟vN^T��Wƺ`��͙���@QHq>E���Uc�S(�l�f-B�'	Mt$� -Hn������q���Y�д��~��\�[8ßz�5Cߏ�VC5�˿2�c���69��17bZ۫k�����6�x�ٺ�K2"r� l�న�"�6�R��XO��2�̰��q��0�{{�= ��!���4�\�>1�rCV0�\)�a��֋}2[&7׸�l6�f���f�i�R}�x��'�i�"�+�OД�EG,�����j��>ni2�4Ϸ|�1f��Ѓ6�Nf�{�Kf���{+FYI�Ro��q���18���wZC5������ݿpXᨚe'�KfX`�;�-�����~ޛ�C4��~e)$bB�
G��Ze�Mv���٦zHØ�V���C��\�40�ky��u5o�;�<2gxc7b���K[��[-�5�p�P�E�}�)e�%;���2�oN�T*��e8��if~~þ����\.\��۫�����΍�!GE��b2��c���=��N�l�}�vn�҇K/���.������8���5ۯ-k��n��q�����<y�v������� u؆�4z\�_nŧ���3�n8lv�qɎ�j�eq<��ȝ�z���Յ9���.m��v��H�+�Rn������6�jCV˜��=�is���Yt���4\mϑ��a��D�u�M];����,$d�Kom���_9���y�3d��#�����]cp���nm�mv9z��qӂ��Ӿ�-�bH��)��f����
5G�o<ni���u�c~ �i���>��"�i�ׂ��p�Ñ��1�ɱ����ÿT���IL�;����0�s�*e-�a�c�4[;$m�%s�s�U$m0de�n�����|��Majq��~�z@ٴ�s�ѦRe��W�S)f��jo<�6�	��#�AcM25�#-1���ͦY��W��4e��e'��x��e�N�_��ݛf��Zs�E�G�l$��+�"�o�_Oi4i��e:�����ٔ6��wע�!��)>�:j�I�i)@�I������w�miGl�Hۍ9��o[{ns�[Y������гi��>�y�>rQV�Gj�0Y�Rq
O������Jg۾w�He4�M�����Gi�m-b�4e�F!�tj��$I��#��0�p}��"�!��Q�n����F}=G�u��T�:�x��;�6�+���92#pB�V���X�b�*'���{�6
�Y2e�bW*~&�q�WhL���{��S�Ղ(�b��E�>��f���l4�f���o�(�-2�?sy�f��Hm-���l�
F�d�����痍��Y�JCx��C�!I�o�qp�2�g;��F��r� ��&�
2�bXi2�`�`�+���RZG���2�I�c[�أ)2�$i7wߺ�y-�J wޭD4p��BXrcMB4�U���&P�S�Fs����M�{���e�ƻ�e��B��S'�ݙw�mqE;8ѹ�Er��[w�7o��wׂ�g�[��ub�2����l�<]���߭�C�L���4��L��/�[%�IHwѣ�	�������ø���Jg�DƼ$P��M�cH�5_}ѫ> 3L�Z���e&P����[�L���n���!�O��s�^}�KIF58�f��@�߁�C�f!�^�k�������`�;^��5Y-(~��r�q�rΞS�j�GMM�\�L��ڪF���ԴZ���������������v�娩6:S��{tD@@F�D1�2�+X���fow��!�})>�|j�H�ZD r��$%2�J@C)&li�M'��L{��si�4�Ϲ}��i��I�����Il�x�=Y�ѦRa�{�Y��dƔ�[�Gu�aH�o���������6�fҐ���P�P� B�ύ֑�ghP��������G+8�S%m�.C�λ[z�������cv�<vڴlhY�T�ex�*?_�~7~��9u��i-�JC���e&P�������i�6��wע�&5U�{<�r&�q	R17N��vu��PC���u\
�,k��V�E߀ �e���)�D$�j���뛼�T*��}>]ᙖ�~Fen�����i!�	�����;=�uK��.�.O����X�}H����W띷�W�L��-��rs���;����>��
Q>��| �[P����ܓ���#ܲj�r��H�tI��2D20b���P��y3�g��{��1M��`�Lfc�{Ỻߨ��e#��sv1�U/�ͮH�@�S�Dq���B�F�g�wg�s�I8w]�)x���d�N�7C$��"�"�0H�	&�7��w�iuܙ��n���x�3&;�.��S^e����@��׻~Ν� 3�"��2�سHe4�N]{�)L�R��0�h E�������H��TEAX���Jg;�i&�I�9�VL��w�Y��(�)2�'��z��e}���!)b2�.;@�^�Rr��0�a�5%���^��\�e'a�r����}i��R�\!FRLMhi�>�H� 3�2|s}�ͦP�=��řC,0���h
��1�QS�ʴ.���jtj���7�8=X�eYy�$^^�B�
�3�4��Ց<M�mTGTD�٘�iM�.�
l���[���:�am%<�D�9z��m�NI�৤ս`�3�tGc����L��v���q//���D�l(�4��e�ָ60��˶��K\�wY�+C�d�.�e��%n�&K��m����e���Z�v�X��[�������ܽ��85�7;[m{����� �{Quv������x���{������ޝ�<n.:�
>5aMYᗲ7n���R���|^>����vO{�����<��Zi
R1I-(
�Dj3������6�vY�Tt<�郠9��{k�[V�,>��k�.j�������&�Ɋ��C	�0�k���sI�4�s�,��	��~;a��0w׊��ha8OIE��[!�JK�#h��]�#¨�"r����44��:
�k���w�+P4>�ƽ �)����,�i�wƬ4�I�0r��� 9B��o����`��{e��h��^����a#jM�B=/��� 2}�s��$����d�<A�w|�A�Eq����e����CM�E"=�;ۭ#}Ta��Z[ﺽ`i��WS�8jL�
������-�Y��PFa���Ìi�!sB{,c�r'C6���g4At/1-���:��rB�Ep��o� �a�B�p��[2���Q��-%'=�����h%�?2��1!i�$,��U����z$�ple�W	���Xfs�Wy�j���\�y�:TF(��Q�n/���W=u[�X��9u�T;Q����"$�l�<�D�ȃOpft��q�*��" I0R(bL"edDb�A|
ec����}�s��&P����fP�=����Q�o�~%�f8��)��C 1����߾;7�P�K���c�#MB>���`ikH���>�\�4���f+4�M'�	i��|��e0�ݿ6ea����Va��
�(��"�����L�`��Ґ7%֑d4W��,�M�� <���6KfҐ�/�FYI�)>��.i2����w���y��t�]��[Ν��ƫ��Kvw!P���q��'�qk\�i�++,�
�*�ɴ-6�O����e�JB�WqFYI�)9�獞�;L���}���ō a���|0��!m�b0�qC`k&�+�SĉI�)9�u��'�i�>���([&��4OB3IHo��5�[�8�-H*;5�Sݙ�E�q����E���Ո�z`p�S��eduݽ�{
2g4R�����/�n�wϢ��5ݹ�ha��-�D�£�u����oT��3Q���&M�*�y�D@I30d�!IF�PEDY���?|{�7���a��i)b�5�X@�.s�Q7"�8@d�H���|[��ٴ-4�Nwƨ4�f�����Q�Re��w���6������[�HXQ� l��V4��i�G�zl%�II�D�g�P�e&�ޕ4�CF���ch2< �=Ey$aJD��"�d��n3�;\ۉ丛X�!m۲�{Ʈ��HPPC��p�%��p�5�)
;^�e&P���<ni)%3�_��Y��l��/��%�IH{��[8Z%Ą9���@���=� 32t��.�����RCW)���N/TA,|�l��>֑.߼ݍ ai�/�[%��ihs�ѦRe
"}އ+H��sجvDB28Se)4���B�|Zs�3A��4���b���(Rsu�74����s��k��7]�^\]�j�Rݗob��O��:��9�Z�����)۔��bJ����C�~���w0VN�8#���H2��a�u�罣��7�n��d�F+"�#P�B��آ�&����X(���k��,�M5迉��LnBF�6�C o��a-��s�*i4��;~l���%��0�;I�l�(L�OBv:@ޫ�g5PtZ&g8m�p��N��6�{N��E0�J@B!��#H����%��+��,�a���[����Éh^+�P�ZMw�G	����c��_`���a��~l�x2|��3�>�r�"���}�Gh�w��%#��eI��p�ds���4�I��+���H�
Ns�*m4��>]�@�A��w
�)�q�$��Xi���HW[��%���7���Z`���Z��hI��7�=l6��2x?2\�4䁰c��tA��;Ҧ�Hi���s��!l0��J`T
� ,z��)*���ElYk���#Z��C�����8=�_����\-��JH{��*�sz\�[�`[�Md䊧����ɦ0o|��橉w}�jF��}ہ�x",�Vmd���j�)��1.�`Ս�N�����R��1o0y!$��T�2�[ՠ��'>�v���f��"zw�1=m��'�p���Y��FgB�՚�dL`}�_��]�q�l��;����m[������n���k�7�<�G�=�g{V�QFj���YT�j�0�(޲3s3^���b�e	p�q9J5ub
ECVpq��cٗ�~��Lʎ��DO����*��v�SE��Q�>SD\��8iRZ��-��d�!�52�NF����#!��;tN�mH��յ�"r��<?a�r�ɷfu��:������[�2�g�&�4��r�f>��%�x�j�����w��R��?[��/�����z��;�b��v .zz���_;�i�h��%��&�-ܨ^�����p�e��&��]巟�������i�tn�J�L�r���*����e3Wu;�<i<��l[5���fv��+̩�~�<�V]�q�Ċ�OR�r�DA�s��"�/���w��6�U�_�`w�G�AY�w�9羹����x�-�/c�f!�7V���]�ۓg"<!���O;�fѦN��<��~�ż��[�TXU �G�l����L�0����m��K*f�iH[1�Q���ɤ�¼U���;�{xg+�g�ɯ�m9H���}��$7�=�Z}�:݆9GTC�?���� _��m3Ck�ؓ��Íxǜ+���gnHbK�I��dsEc���'i,Yy�:)Y1=�G�A�X���w2�n�G7E�\�(rق��n��y��B<6-lj+�����s�]q��ݐ��ݺ�7b8.f�j�WnKW7'<N�>V:s���V�v!벞�Pv��Es��1z:{v�@;c0[k\�l��9H�&�qv���!\�'!�{�9����:��&�!B��m���a'v��X)E�n�Eú��gp�6�獖싎���ݲ1{mѦk���C`�ǋ���.���瞱�"'k:�=XB5ڝ7wn�H{q���2g��v�]��Aj��v*�ꡕN�k�:7���;Zk$uîƳܺ�n{q����%i�C��2�����e�u�{Wsn�2\<�y��Z�h�H`��l3�w&z�G$�V)��5Ԗ|Og&�F�q'F�C۳ў�b�p��ی�#�^<����e*s�;�!��X��=��P2������`�q�s��p��τ�쩚7�[pG���-s�{Fz8ǘl]\���6�����n�<n5�m���Gp�!N9�n�9���ūX7i�`���ۘ�88x���[Qq�V��u�Ks����գUq���#�F=r����K�l��D����q`6�O\��ݽBx:���9��C�+f:8�ݸۥ�Evs��1�[�mFn�p.��7Xį��l�^��$]�dw�oF����ۮvKg+ug�vuvEq�k<�f$%nŨ�m���,��cK�<�����v;X����"@r�Е�i��m=�h!���t���鶺;u��5�./`�/]1�\�q���W;t����8�ֽq�Lpv��� �z�fU�Qpcmu�Nˎ���ə�a��c��h\�p�jut�ݶ耗�=�=F�ɧq��\�Y��h�F�X���K�P���M��G�.4��p[s����7=g��v���8��N�$Us�Ӭ��n��\O����ݓx�(�+w;Oc]�y�N��͵e7<6qQ����vc���Iq���n�݌���'��:ĀY1.kc�J7�X��(�NB7`�:�� ��x�׻./��5������p�vT�gP@Ӽ�Z��/7�l~n�{ 혜C�:�Q��TJ�P��F�-#R�M���HFpvx��2bC����a�-�Ll�yfn�f�l=�,>�O����=�F]8�Vtn��2�F�u$N�nP*���h@��0��ɲ/�n�$���.��/v�����2����_E"�������kQߢ����Q��Xɾ�� �Y 9 ,ʇO\c93�X{�~ْ!�z��:���3e��v]�$�SŖ�}	h�2�l�}:�gLX$��Lh}V�$�J��b6����94S�2�`����\{la�9ֵ���ûv�Gl׎Z.HL�Ҹ�$�z捌IV���k�>G=�ã�;��V�a>;'v^�@�=;8#sFnB�8~�7	�l!��	sl�P��Fj'
W&K�HE�P�TY:�|�
�bi�+w����k�l�@�dʣ����:p�IqΚw&���U�M�m��^���C_?g��'����~^�2I�ާf��bK20�q �n�jبԄ���j��[�0E���C��`)�~(k��5�W�Z��n~��X���ߓ�^k��:�/V�Z&6���l�gu�tW:v|ŀ:D�Lu;�Kp�9��������mѼ��َ��
����h<vL�/ck��r���nCZ�Q[;�zT^��N��q�$mq��n�&7���Y��#�d�{F�NҜ�Zۆѹ�]t.�q0t>p*��I��8��r��3�;�q�O''l)U���n:�����Q�s⻧��1Z.�{"�b�m��n�ݷ�2�)}u��LB�I$�a���{���}p\��3�pnE�������sX���X;Kqq��>�t�Zu&Fٷk�&�o�e-#���]�&u{x�i5��㶴x�)2�'9ε4�CL1���q�W��n7(F��,�do> ��  jR��
���s�ni-0y^��@�
4�F�j2Ҁ��m�a���o��0��{��M3�A�=�p��@���ȻHy"�qX�8��~�&S�Rc���m2��=�}����gW����i;W���(2,��\�z�NIQ:��n��CL��,�a�Џ������k�*KC	���\�e0�s�1��b']���ݦ���v���s[�.���������k���m^�=E�,��H[&�}�ņ�i0���Z���o{�= �0��<�Y�2�	�����b"�(�ZLKM!�ӬJ�&�>��^��8���yg���ʧ|�m�����R��Q�U��[���uZ}gn�N��t�<�v���j��6���4D����^�]/�� � ILXD�&a�i/;�˛��&��gw&Fߋ��r�]����|M&P���Z�	�^��gSi� k�B}�t"���.$ a�M�da���ni2��;�rY�2� �'����&����	�0�kj��`�d�L@Ғ�H����=��#[�w��L4�Cx��C	l�#I�s�n�F�������%I�ca��:f�,2�OM�3�&��}�{�C,w�Z��i�\=1��1N�v^{V��痍���3f�[ر��U�g��a��k7D�[Pt5�#�X��w�{��ֵ%��}�����\�l��_��w��j��b)��RJV�(|�{|퇈P�����ou��Xe��5�Z�<I_B�]�Up�hdBܐ�i@�@��`��4�������/�w���Jol��ү`��t��6��;����z���6t���t��3��S��Bg���{_���;�yk~�⛣� �%�"`dH"�
K,�����@"O{�#@���z��ǿ]{�����0���]��IH�"�RF��e��	I�{^K��acֵ_���{��L�I�>�}�Y�'��ħmƐp��]iZ�BPd[0���[�nm2Ͱy�f̳,0��s�]i��3^��>�A����e�oi�"F�0;��j�F����nև��y۶�;�u��`�i�d�'(24�!w����4��;�̳,0��{����Jk�<��ȳL���c��2�Q��4�f�8�=�2� &�Rs�ג�L4�C�R�JC	���w@����|���	��#q�@�U�w�.�7���B9H�|��&X�;�Y�#�����Z��ba�!@g�@)
�C	I�g.e2����e|��w�����wɬ��\MtQ�|Õc�e��;;�"��b�T��T���W�����ɼQ\��&�`lLe���o���>�b��Q`��
�R��-FD�IF��Pd]���i#F�4j1��w���r��CHg��e��T�&��ӈ]F[ϻ��Mz��S���c��g�� i��	a��*��jD0�P��P'�gM��ٺ���v��M4L�s%��ٕ������6��$�A���r�Ϗ}���f�'{���0�a�w�@I�)>��ۭ#h}�fT�1iI�c2�	��;�a���Rz��RO������a���eHg�Ro��x8 ��
1��R��CHd���%���Z�.wf!l罋4�Xa��"@�K;�(�`��$�A��X�]��L��;~l�a����Va��%|���%�u�Ŏ�
S���,���Ex�(P<�s�O���q%$ֵ��e>`'�|={��X�5F��"2k�1brs~��N�h�P�������I���	�=%iB~���6w*��
��k�tE25u�|�#����M�V�([/]��7s�%��ޖ�Nmv]IpS<%n[��Nv�Й� �>v�+�ٮۨnQ���U�������q�ݣ/L3`��(VZ��'\�1vU�DC��2b;q�y�cL�gp��.��{f�e��q��f���g�\S�1���ݲ��6�0���׮6�{n�=(X������p>M��w]��!�:����P��3�{�ν���6�ш35A6L!�",��c(Z2Ѣ�ъ6�,�"����3�ƭr7
<�\����b�A�7$C���+�]��ܱ��2	t��T'�O�0>M{�sp2�!��چФ�5�Y��e�q�}E�l0�+���P��R���C /�.� BZ������4��o͙C,0��zv��=B�p�@__|���e)	*$�a2���}sIhi����-~!���{�h6�,�8��ZЎ|h��g0��.v�lx��x�!w�ua��4����Y��W�9�카�C4߽�28ሰԎ6�T#25���i-�C���8-��	��*�ZC4�;�b��4����AizRq8��>�9�l�;[���p��k����붡���Ӌa�T�訷��������s�}�9���ti�yA�� 0�5dq���f��@���"�8�i)"��e�ފuq����#�G��37Sb}����e��=k"ovh��cS�C� ��9w0�9��r�ǃ�q}���od���9�/�!L"a����*�j�5DQ�,b�-%E����1TX��$ RE�=�Vo>s�2�k�t͙KfR�ՕϨ�=�4����r ��)�H.��@�!�\��eL��X����Ii���9���&^�B��o7�a$�I6��Sn.����I��7sM�ƕW�m
U�|N������Bj�	&Ȩ���3� ww�f�z}G��3$��흎�S��BSi�c���e�v���㍺�um�����u����e���CN*��#���~�ܽB�,yƪ���E{o�31�;r���EH^^v}�9ꮚ�埯��ic��^�����ވw�i"�Ap�Dӥ��]ݬ:&W�\��L�/@��N3y�7x�A��˥Vժ�}ݹWQ�u7�a��¡]�eç&�����s�B�ϧgc_U��[�!7u�8�1�����4��`�,"�lj6
�(��m�m�h�mh���`�^�o����ϳ�w6}܄v���e2��^����Y��]B�,��5U��7�]�^�Aj3���	7p�zMs� ��fV8}�j�+wT������j��$��j0IPJM�	�t5��6��p"cl"���;.�uΤ�ݟg�<^z���Q��UW�"d��>��fĸ����y&�,��,�[��P�����w�:�W�u
T�Ӥ�{ﾷ�z#��&�&.i,Z$̫��tkG�>���P��˔�^��fPKAd�|����~�j�zx��W�B��u����bhg���_�Y��p��y�>��&"��U\�O'B��F���wsj�suv���6m1xon�|���~��M��@"�m��U�ѣ#n\أTl[PkD�j*�}Ó��4Ȳ+��`,�hdE2]ba&���,�M3��Q)�L3{:���+�`��!�k����yB@���Pyb�ݡn��y:�(+������r��&�ms[.�����3h�%:C�߭��i��}���e0����	i1�m���Q�!w��E�"��!}�+��m��1�Rb����ڃ���"��"L�=}J"��#y�+�U���@������M�M%!4�#H���ܺ��s���P�����]���j4��)�Ϯ����J.e-�%3~�~��$�0��rQ2̦�g�3	L�#+Zۚ���L3��r6�R4"8౤V�d.O���e0��~�L�i'~�r\�ZL3^����4��:�>2^^{uu����]��p����+7�r�C��*5-D��#v![ܬ�vj�/�G9��_k���咲82���S�Ҷ�e��q� @��N��&����������8�nݎ�*�5=�4t[+��K�ܚ���ۃ�a
Ŋ�:lr�2<ktg��D�h�Qų�G3��n9�;�=��7k��vuv�j9��n�����k��Z�
�v.���ݍ�$!����=A{���7���|�{+�g���u�g��4�k�[:�q��w`��M��Ҙ��X�Eϫ�ŧ�F��j㆐�ٞm�X�F��F���c%jlTEF�lF�j40Ԛ��v��﯄���Ƣ\�/d����p�핇]�d�;�5�79lQl�����Z"��c¬���i������S	0���g�7�6�O�]���Y�h�@�jy��ґH�DQKi�O}�d���G(V���։�a9��,�(�f��#Y��D��)"uP�sH3��Xg���ΖKO���Es��4��w�.���}�{�"n$a(��q� a�!�ϻ�+Mazl�ٽ:��@�!����h�2ϓ��$8��f&���Y�"��u]�4���>�}��>f�]�1`e�&���2�^����>F���i��R�R6�[I�*Lm�s6"�W�����μ��B�'�&!l`�L�����ܺ��w�wE�I�a>�s��='S��=�}�4�I�$�Bc���1i�t!�o���Ƒ�n7=� �e�P�	߽�S�o�v���ӝ\������m@�=?1��S8�.���{�N����#�m�2v_�~/��ؤ�ZR$����f�X�E)X1�W��^��-��oO�0��g:n]U Цk�tu���܍$�I�4�Lc�>�y�!�w�z��,&�G���e�~"���}&u$#pB�V
�}M�����\al�{�u$���=�4�I�F}����5�{��"�IAM2�i��Q�ݱt,�G�o��f�m����j��g|p[`�
|�)�a�p�2�$�F�&�b�G>^��In��h<�Kqs��6ra{:��R�Q3&PF�5�wޱ�����t,�L�z���&�`����o���pT�����; a�{ϗn�� p�θ)�w�<��Y�s��x4����S���	�1���@o�{�"�sdO�c���^���p]�5 ̝�n����f�c�k.���՛sҶk2R���#j�c����%_)Z�q��iQ/n���Y�w*q�]U|���m���yʼuuÝ��/14��؊K��/���������i����+�d��KP�<���a�#�lj���?Qr��I�N�nU���o�v�BcJ���W5*�"w�y�=}{�@�jуݹ��^���������e�5L��-E}Cu8���T��F�-1">%�m���ˆI�c6����cs1]��Li�=�T�5���Q�i�5���9�&ț�1I�9Ni���vŬ���v��b� �7�n���i�o/��W�QK�{MՋ���E�]��=��Ť}j��o����^}��
����k�R����|a�o�r3��������������]�u����6�PM�C,3�ke��z���f�y�����/?�q����|�{5����X�Ʀ�#<������[�ZL�m~o	#�s`6�ݩ;���j�}��;��ʋa�v�B-�%���n����_6d��<�����'�䚓��D]O�����˫z=�琞�rm�� �����rS�D[M"j�V��᭘3X�%�6���f��Rv.���yt��_�(�jX9�5��zH��O0<�8]�<��9!7�gb��S!��}Z��i~���
4�VȒ�,���a;m��f��LZ5܄p;w������Ke�-���
���E�C��V�m����J�v��{�Q/��j��o���_�5R�G+oX��krQ�F�=�t��]����2�*R[aň#!�W9H2�oX�g۾�	AF�;o����6�c��uF�Tt-d�k�݁�g�D��1���r��R��g-ZC'$ڇ)������p�P,9��6y�1	�f�
u_�O^��^�b����7	h��=������m=wt���u�r����V�V���h��{�C��|$Y�m��wps��"��g����'ެ��Oz���x�"��7��,�����A��,+V��Z��7W^0�^�V���ăN��}�]ߧףoл���˴��43F=�B�=+'������4 \t8L6��K�y]~�0z�bk*���q��ygZ �M!��!��>��4.�}�	��M�ǻ& �l���=1i�vy�C|s�6��i��i�K��w<ՠU�fN9��u�{�[�Ed�fé�qv�*������}!����(�0����M�d�����x��j}���o����gk��#�]|�~���oso�Z�f
�>S���ݙF��͕j�e^��GP�9=��{{�8�C����8�UAgst�P�I�͋(�|� ���SK4����zm7�J��
����{X]굿>�����t$m��7�-�op~�x973E�Q��I8�dH�n1�8L�9�tWF�J+UD�Q�-�cl�`ƍ�P�F�#Dh(
=^;�YĚ`��w���;�t>�d���"��j�T4�J����\��o��ɖ�ΖK|� C^��j��>�,1	��jH[��5�o���4�������|�����R��t�|*�~�>~i�lr�ŉ�.Kv�|C���ɣV�{h��p��i��ra�N�(F�8j�>~�W$�z�/z�,�	�s���o������D�	9�Vs���C�00�����e>I�{���M&��+�~�d�@� �	���kɥ�F�]�44�>טּZO��o�Śa�q���������t�f��Gy9r���C%�� &����i4��=��%���;�E����~��^�==pȑ�mK���T*�Ù�錸�ګ��&��vCS�����2���WA��=[5i�Ʉ9�����~���)?������ɒ+�I"lAh�6�P=O�<n��H���'��b*���n;4�L���[��A5θ2�)>��7.�"��o�zƑZhx
��{���2���sɓ^�� %j�f��۪�]7-o^Ѭx��Kb��*�[7�GBU��-��{�=�4�I���-'��9���U!\�y����}悌�.$ a3wgtt�}�4��޻��ރ2Otwu��do��!����=�ƪ���'����v����k��ȷ��܅�[)���
=��Yi{�����t��}�}��o����CR8DR:�F.�Ͼw�0m8���z����fI��|.TÎ��tUMשq1�L"^Ҿ��늱'��+�����븈�3j��f���WY�j�Pd	s�,�9��0�����o�o�;�lmC��X)�-��FC	��s��WV6��'8��a���T�x���6�K������'hN6e�K����<�����M��\�1�Iq�^��綗Z^���c�ٕwC��ŷ�x�v��j;
3�7����NO]//3'5�l�]+�����w:�d��r�q��yn1��\%�ۨ;#�[v�ۑ�n��2�K���Tm�hط=z{�x��}��n�޴R�c�ѡ(Cb))�D��(A��uw���s�������p=�y�����Avd�s��i[ctimu�z{Rۊ�ʁz�����pd��q������ RW�xUTgp�
H$hEr\߽��Uh��}���{�wwy� �*E�[L�j���31[�'�����3;ު��PxAL$�a"�m�π��z��ސ�;����(��ye�{����ԑFS���~���< ����{�fc��uW��Q�� ;�Ѧ�dm�<X��XA��t6��{kj��n2��	k<���q��]�߯���EP��31���3�u�nw��M�Sm6I4����J�-٬��u�0�g�ǂ��k��y�pL�#��y�%�
)�=w�Z�{��j�o��E�Tw	�3�{��7��l��T�+���/w�q�Z�:�Tb�De2H�$b@(�1'�����}�����>�5��eW�1�l&�Yg�xHwG9/�(����{�fb�drG�%�l�d"�U^|3ޑ1Y��T=��g�|o}�S{Ϝ�I�W�Ap������ ��x��{}�Y�v|*�~��H�4[eI#	��gqh��=�ݱ���
��0�ཱུs����halEP8YN�w�Wg9ދ��|_�kw�w3����%�1�������y����+7z*���}�s��DÆb$0�lUGw�8����wyfS�Ga5a�^̨�c{�۩�i
�ar6u�;n ���Q>�|���"��O�*˦jnwK";fj�5[���ź3�Wz�s&@QH�FAAH���X�@g;�}�}����sD8�B$C
�����s^��j�޾3��ޅrcۢ
�R`�!H��s/��9��U_O��7W~���w����E��ZM:%��-'��,Jѝ�2��)���qP���q�ʱ���Q��v6��6�-��w��nf��E�~�}wϺ&b�o[��"����E�lL�{�5Qz�G��I���im�C,�������L�}�ŝ�u�6k1� �*��I�ӊ�߀��x���~2Nf��vK��=]�:�
2�'������5��Bb���!����b�me�0y\�3n�&i_Ě���tDSb������8S٫���P��@
5�|5�Ȋ��\�G��g�]�)��,�-��T�k�y]���
�Q��5���j����H���Hn���ɹF�b�*��7O��#�<��n1s]bh����T�j�4Oo��?���)���4/4O���b��*����A��Pa�,U�ފ����x�I��d�ͅ���뷻̂�(�R�#7�̓Y�N�/gP�1������I�栂�4�M����,}�jI��S&+=�5��f��!�s��M��Ъ>Α2|>��蹿x�ʪM��'�ә���>����^D�(�8��7w9znsL��
�xu��ʨ�*�j��9Ҧ/����������CџX�4��+p�S[�p�`ڲ6&*�N��im�����p��33�̡���5�Gk��[���]���B� u�s�Y�m�G��m<����9�y�ktz����U6V�cv�&詏b���ջ�r����-[�<�,t��GY��5�n�et�ն���X�l�u��v�i۴ⳙ+�qh�@͸�a���K�2]��/k�M��-�ݬ�1�ѹ��7�;g����sunƬ����g�V���ח��z�⫤h$(����fh���_?��n�ڞ2�Z�8��#ю���8�j�0�����uܻuի���\���g����U�阾�=�|.�o�L��:a�����I×���^g�V>z��_}����s����W��j��@�c�s-��U�>�J7w����URszy���r��2N������t/�ª� ��.�o	P��XD�Tcsx�׾��yq�ܜ����r�U/w�?��{�ߡĦ�X��ɵ�=:�v���n�\Jv��Is^
l�h4�k���pb��͌�xUQ��z*�����}T�sx�ׇ���)�me�U7��������=��W܈��9U��n�eE��3�W!��.�fK�c���D:��:����6�z��_B'�/��P��}�b��kW���y�}���*�X�F��Q�c5�dFU���8��ڳ<���ox��`�`�)И��E��z��t�;ДM��Zi2�d2ʅ8���w9��f��=�����m���)�9�������F^�qw�w���I��a �L��)C�����i7[A;y���on� ��۩]cJ��7$Q`�Ql�Ǯ�-���;�"d�^i��no�W_�-/}�ׁ�2�1�q���'pw?}�Q�ީ���Ug;����{��a�L"ۄ�������꩜�`���ɕOb1NA$(UP(Ju�9W{F|��ә��gۗj4�]}����豢'x�+�P��v-��P0vF��?t����F��)]~ dZ-QlW�u��nj�ET\���-�lj+Q @&��_A�|�ï1s�z�-�$m�,$�n���}�1~�yUooH����{�]�2�(M0AF%�N�w����y�U����U��4}������{�u���������8ç]פ�Z.^.Z�;��ι�-)WL#O����ޡ^�p��UM,;޿|>��m5Y��䉈�lG����������7-k^��{�O��
[� WC����p�L�����tcy�|����.�oz�M-��t�Q��fA�{� �\��ً{�*�B�Ҫk�Myק_�׹���8�pQq���vV�t]U��fVc؁(�y�EW����t>�\���`�j~��ԱH�ZW)��y-�g@����6y�S���]��|�� �YIUk�卨�*����,����("�����X�=Y����\!�Js1k��ט�B�}�To�*�����:\>��p'͐\|K����A��+��,��lm�wу��]=x님�+y9� ��Aa��^��U4������߇�J�[��Q�t�^`��m� �LS��*�>�U��܅:[ޡUJf�Ί6�?rHT���6���v�����}�ǧ�b�(�xUM(���[��"��u�|ޯE�([�
���{���>~�v���z�R8$q�aɷk��:^��{|.��5Ǣ�,��URa�o�Lq)���]�����u�����q��������n�vÎ�^�n�*��V�����5"�)e��HP����j}����uZ��ݾ��E֢�m���6jTs��WH��rv�i�A����=�ۋ7�~�}1z};W���EA�Қ��Q��bS������Ƌj�_y[f:n�p�j)�rd�;7��w�<&&��4�'�jWۊ��w�;�����5�~Z���(3X���(p�A�g��y]sS��>�몫l��-�.�����d�9\��Tn=M�_\�ӥ�������tU�Սu;=F�;ı�C�Xi�⨾���Q4e��u�m�{��#�_}����އ%\���]sS�Vwf�~p�6��@��^�c�i/Y�7�o�k}��r|�����!��kN�y�\o�s�3�fc#o�ۻJ�Q"���'f�P"A�{��U�֓4�E�_{�_���;���� /�!��yC��m�ziD��<Z�2�B�j!��9�C�d�ա{��uހ`�g��B�`���ٛ��x��ŉ动n�Hͽ����5$�)V��9����K�o�@���`�N���+/kbj�e��a#J�א9ƨ����l��/��zV���rM�u���؆w�"�5����$;�<����Tyi֜U��x��c��+]�w���q�����2#���_ފ%�a�n����k���$f��`JW�[�S�^��=�'Y��d��^[�΍Yܬc�mw�@}{o�D^tn�>P����E�?��B����{=�q�-��Î5�6="�äzsvo�Q�#���E��������后�i��l=�9ã<A<�b����_n_�f����|���pBԐ����O])�w6���<�׷<���g8ۮv��B�y3ד�S��0�w<6�W����gG��
Ev���q���vL��u�2�㵴d�7\p��OrvP˶:5�4F{�ua�tNdN	rs��e�����Wz����8����%���S�uU����=���6r�&��`��3�n^�3\v�v��◷\���6�D�x�Ƿ��X�7zB�����m��7�Goe�v���U��&,�rڂ�ݺ�Ф ��'�ivݜ�.�����<��	�M����ͱ��v����Of8�rsv狜z�s�Ѻ`�td���3'c�n3�v�FL�	ˡ��1,��h���.4Ԛ磭���*�1ϞS�]�Yǳf��u������F�XH7C�[l�Ħ�7u��Ewvݽ��n�݄�槽�נ��ǥ����xm�{v�`��T'uر�7e���=vol�v�ĜX#��#���m�s�rojҏ�&;� .�wf�؜�mD"��]�/4���u�ق�|m9^L��l�=>�W8P��\�gq�69�I����2u��LO��ㄎ�\�[��g�FX{n��Wn��ev���f}�#����t���3�8u�^����dw/���O�uk�ö^؝�=��i5pl蹺3�Mw;���q��y���rS̺]�vx�u�k��%e�K��7	�QA�s�1�c���[�c���ȕ��� \���5�<`c�ϋ���9'�ɸ}��k�=��j������-r˥�<$�t@�`9��与��m�^�p6�=�4s�F�.�9��֫Gu�=;�����O']��u�^֮4��;���{V���t4m<>N�^����qtDIk�M[�n�m�̏b��v�;����e�-��s�s·��e������e�Kݝ�^g���R��(u�c���Yx�۞�P27�z�n��p�e.:��Q��{*��1h��KQ�l�;&64�Xh�[��eݓ�Bm�������pn;1�֮��A瞪�x�����l��/A'4�Z4���i3���Ѭx!i�W���]?W���	.���,b�#VX���7JT9ڄr��F��Y���������+ٯ���ٜ7u�|��0�\CZL��'r�ʿ	��w�ۘ���Y˸�@�u�CAX�ծ6Ǽs��e�����8���u��e����r��4��r�A���\zz���lQ\p!���;4
ӻM���3y���!���2~�D���G`�z��vOal��ܽt����h�P�3�� 8	~Y5�n$��$�|=�x�"��MoX"�U+��>�S0P����y�to8c�&V̧y{�D�W�Q4���%s~�,-��ŏ�yz�ԓ��_��W��w�$1��LL�tԁ>-�|"����䴎<({�w���-M��"�K�N��/<������O�����gv�l�`��H���NW��Ӵ�l�`�^��޿_\|�&��a{�b��cN�?�ʵ!뾬#��	`����!���⠶��b��?���'�M�7�M�^o��tqUP<��y��</0/v�za�X{�)&�*�EΫ���y�>_%o��u��C�٣Bk2;����*Y�r�>;�@=�#zQ����+�L+��C;�<}ǾjG9	<2�,%����/���2���bf5�7~�N��"��;UWhq�x�;�.��O'�O��d�s�N{RJ���뎶2�Ɏ���ےγy�eڶRm��ώ�;7gp��u�nċ�m�.3�����:֘�q�%���<ޏ\�5K���\�8y�Nv@oe�7�+�����L��m�9��Onǋu8��*��tۓnQ;	Ľ��-����1�v���z���[l�{W��ȟ��TV�b�b�E�5�cX֍�m���ҝ�!�Q��l�C]��� � z�������x�f��6� ��ԎMA�i8^�[��wkL�K0n���ǧ�B�[��P| �(�S(�Z�iD��	��]T�n�M-�r������|!��'	��&It�.��;�Xw�S��n;|.�<z%�Y~�A
0�$�$1����|^�3߽绚��v��>��k_z\BA�A�)�)ҍ�SK�����i�Ϣ��-�B���|<~���_��g`�ySwWl�A�q�[Y��!�nu۷�7n^�ڶ�7Eg�����n�5[Y��O�T��5UR������ed��ªiwx8��	���,��qN�l�+�P�b�c��N^om�\�f2$�-�����f۹
�h�)oe��&|�&T�An�ގ0��`j��s�����:����1{������72AH,��li+�Œ�Q�( � � {�q���o8{�w�k6���� ���F�m���CWv���S��*��}���Ǣ�-��UR��,�A�p��//;T"�}��f���۶������T���6c�_��h@��A�[sk��N���oW���-ޅSJ7�un� ���E`r�m8ʐ�"l\��G[;�k�v�)�]g��4n��я@��AA	d�C���׭���3�}�&3�p�}𺷍w!N���D���4�v�n�*����g{�.�i�R�`՝�a��
}I����a'Lg�xeM+ku
}��|�z=[q�]�1�◕����a�{Y�{�t	j��ET�\z]	٨pg;")i�ZF�,��ݨBou}���<�;_s�0�d��E$[TkF�Eb�klh��� 	�>��,fc/y�����w���ۍ�-8�ٻ�� g|%3�9L���
���������&���0T$�:���~�5�s�o[��r�}*�B��az#X����b#g6Ƀ�������	P+u�k����RD���v�Z����<����7ޯM���8̾���+{��s�A�T#�H6�q5{�3��;9n`�>�l�{���AL$Q`�i4Z3;�3y���ދ��������ڄ�$�E8&��|���z�npy5}d�ɿ{fm��>陠���Q�U�X��1�r,c��M.�ۢ�S�Ӎ8�^u���ti��UӮ�������_^A��kX�F��#Tm�� �E�AB����Ƶz�o����L�����������)s���3��\��7]ݮ��?w�FXm� �Oe�4��u�m��]�yuĝ8-k��*��d��Bm�-��p�
i�x���UM+ku
t�P�>��-ޅSKw��T	�	��ٻ�Q�3��M��s����B�(��U��ow��L��p�h2�)�)��H��
�
��>��x�U��L�U��e�l��H�$��� �ޱn�n�UM+kN�:���B�Vn�0!�BpNI�SJϽ��m{���U:K{�;�Xv}�6�b7.]�k��Zz�^�hZ��
o\;sQ�����_X��u��5鎐���p��ڊ޼p� )kwc�"^͍1%�G<�@m(�ƞ��A-�#�q8�u����uq��q]�f�Ƴ�>��˻�s�@`9���u�Oh�u���:;)]]��U����ݵtM���1�E��{6�am��e�Q�ص�:������N�>�ֹ]܎�s^��t��l���&G���={E��v��m����w*���vs��\{��l�>��,�xT�n�E��g<��欦�[y�����F�'�lݱе=�;���Z,h��5��-b�`5����Ο��Ź�
���V\5�b{@s����0Z��rp��b.�εZr��:u�S�%w�����r��)�ޑ3*^�}�ռ>�������ȅ���%n��xy߀1��X�J7|*����b����Ѿ�+�@P�h�wj����g�����8�
�)opUT��	+YL2ڂ	B
b�p�3��X_GE:[�����2�4��Q�A��[�3�'��<軖�(	�z�/��&3�x�^?UW���dA�>gu�؎۪�݊ZN���\@]�q�Ы���a.6#�	�6`L�aٯ��wj^SJ�����X�|&\��!�i��%�,��������}O���+<��ݨ���v��p<3�S\n$L����<�L�Q׃ȩ�)_9�2;��È
��>���Lҹ8ͫU�x_N��`&� ��B,�� M 4T+7|^�Ǫ||rgg}�.�fC7�>I-!lI���矼���g	�����rp�)1Y�: ���P�䉵�=T��Ⱦ�"�59|��gz�b<�}d�N6�8R
Y9����ֳh*1�ܪj�^ĳ����a��7*ㅦA�YhJF@����Zڬv��Ý�g��nx�q;�Z�+�9�]1�((]�9�S�X�U:���2�n�2m�Rۍ� P'[<�u�}T����K}�T�^i��
���P"؃CJj�O��fI�Хɛ1y�������ħ_YPTr�H終�_l`M\�j�͞Ҿҡ���wz�p9�'�'W{�����;X��\��%=�gxq��H���dR@XQ4H�Qso����3�w��C��,�ۊ��-��T���55z}ʪ|*���̵�w�*��RQ����ݩ�}�ѝ�7tw}>����&O�����4IA:ݲ>�;;@t7<,y1t��:졯%�e���鶋���OgGjGG\�??~\}�U'��̓��{���^{�iv��@,�e(�
��w5�v�s��U���EܨY�UM,>�U� *��3q
d"!8�J�%��UT��Ч��n3��&�w�3��Z$��L2Љ�3=T)�>9��T���i�C�G��K$\�Ӌ����p(E�ٹt-ݽ�����ҍ1��G^q]z����(ın�M���}�Ǘ����?E��5�9�+��`������A��������l��bA)����SG�����z��Ǽ�<�ڪ�Ǧ��I�(�T=I��N�V8�iN�$C&��_�}=��e�z�����Kd�h"�P�MCI�SX���4��2k���Q����!����$��N��P�| �p�x��Y��Ws����T/&�GA�Gr%Q0��ǧޱN�g{������-��z�U(W�hA�T#�Pmʩ�
���O��f�s��r�n�U\>���X�J3��p�MAd��I�wV��P�K��B��,ͅSJ�w��ڌ��읲a�	����;�4.r{.V�9.>��fd��'�0���z��DsXKޝ8�|�
�k�39���U��̃��ӹ�/����۹#}�ߝ'ԷV��fs���mbr[�������/��7���{W+�b;n��݋niێ��z�7(�b�IΝ��͊)�����,�dӮֹ�ʼ�2���؊n���v��z������ol<V�	���3�a�Y;]��竌s�sk��Kヅ�b�����]���E�LK�x�w�����n�i�"�;^6f��ܾ	��9���9�r��Dn4N�v������ۻoeQ�cF
�n����/;��w	M�;s�]���d:��"�8㶴���]�]�u�v���y��@ʶF����/���U+;�)ҋ��o������B�%�xx&IGq7u���/<*�g˾{-oE�\狾гU�o�v�)��h@�L�*�f��M=�)�ﾷ�B�T,ͅSK��=�BqH[0XQ���
/��䴷zU+>���{{�3/��Z-7��h3&اKzḒ�|��W6���Tҋz"\�����L�� �9�a�\�;��s�竍<z��M�=�,]us�5W�-�.���$�3�z�:Q����֞��� �ɞ�3+7DTI�*!�P�%8U4���S�Sޱ���&��srv�3{�����H�OS���Ln��[�^B_��u�?v��Y�����L#r-ɩ���l�9��X�G�2nlۮ���cz������(1Ub�,��$D����^1�o�q��̙𪽜�����QP��|�o'��
t�dL�ﾧ3a\���USK3Y2�DBpD��S����򻥇z�:Q��Wu~�ޱn��޸&G����c3.�B����j���ڌ�2�,�*�} (}Z/Ĉ���i�M&̷�뎂sq�����x��`�3���sg�G�Yf^����!&-ڎ�򻳇�B�����v�B�7�8�耒m�%"�������)[�ʪ��*Tfg+���>)���-�T-�2c�}�d<�|V�`cļ�����3�g��M���=��*�3��͵�+v�b�ubbvƍ˷"���0 Z��y ���1R/l�V�KN�-̃��0����xL�q4$�J�g/�{#���.�����p�n߈!ID��^wے_3y�Fc�6��f�v�Tkr�lSr���Qzr�^�q�B>orY�t�{��/7����~�������m�'m,���V���q�/=�Vt���๞��Ah��.M�L�Q�f�"��w���H�4_5�2��̵�/�lmy�<�Z5���P��=3)���pv�*�b{�_Gw;�<�˞��89�����jd�,��3p�u�xd�ܽg-y��q���i��QL\M/����;<>�&�՗S��a9�`�O���I7$���ĻưѬ�髽��N��p�����M+c2`٘�7V޷�(R�!���=�ã��ʥ��i`5uϱV���&��Q���=Om�䜣��H�Q�$bFN��ާ�K�:h���th+ ɧUc��l)4Vd�[=��='��.��p�O�����9������3��_������m7V��i�×&�ˢ��Ԯ��sW��4o��}�}<!>Xi���,�$e7������۾����r��׆Z4�}^ٓ�z`�ѵ{�q��i�*X͋?	{߇H]�qA���qNm���1�u�@�=�xB�_ªE�d��z��=�KYP�*-Ol�W r+�H1����\�CT:��1��i^�Sktff�ˤr�z��C^�'���a��씜>��>,�'��p�g�����@���}���K�<�䗽���I�OB�w�S�Ȁ�N�AC��]�� ����2��?2�����<���L}�Q��ϓ�:"5����/<~�R�����ත!U�-�$a�����^��m���C×{|�����'3���$YI�Z�Ե�ظ�X��n�|�SWg��ۑk�[{��x��%��2��FN�w4��i7�r�h$�kF��jJ����&vP{�-gqX0
 +F>�����X�Ui���,L�[e,$[!j*ˍT�'EGw����Q�-�p�������6�S[��	�7m�kS
c�i��fh�^�)�pт��ڽf,���޽.�ʽ��լ.�WТ��'D����o<Ƙ�,ؚ�]5u�&?i�C<��9}��!�x}�qmTcn�ę�}�,�ۋ������i�r���Ky���*�-�s�T-:c�3�@n�T\�}��q7��M����\���� E��AAǷ[�����XQ!�0cеizH�8g�gMTvd������(ݤM1H����x�e�l�xA�tK����)�����4f�>��cxx6	9qy���Β�+�S��3�����7{�=����㍧�Ꞙ�s�'.p�Pe�� ��ӛ����v'��Ü�Ͳ����gDx7�m��0�%�`c�f`��VRqkZ�Q �Zy�3�8�~#.5�Ng���Sh�"ȌT�IEǺ�բL�=�F�p�`��1�sw��OP�k���]�^O��w��~^�JT+�4 �*e�Pl����G�b\�{��]���|����T�����?W�i�������]K�F;Y���Krp�[ebz<�/N��;�g,"mFec~S�n�����d�����M珢�K8.Bl��I�)�B5Kw}~�}����U:q�֢����+���~>��0H�8��&1�a���f�ƺ�����.g�T������Kd��q�p) ݛ�*׽�|\͓���6n�=UN�O+��A�:d�*�;�m�(☋���1�rz��=t6v-Y���a��UCdV:P����(t�ՄfQ��j�����n��5��}�s��E"�E@�&�GV������#}��Q��Aʳv�.������Y��OP�t�wiY���|�x�,&Y�F@�Y�&ջ+��-�pv�e�h�,��]vޗ�1n&�]��,�!�	 �CH�F<���N�<ͅ{���/UP�۾>�Ǐ>�N�T4�2��0�ݬ;"x�>s=�.�x�x������
{w���F�0�bi8]�[G��\�kD��T�#��wP�������!�*܏�j��Ӿ���zD�T�6���|���99��ࡘp�BpFb������b��w>T�����n��Nz�Y��v�g�!�*���q�3�ǌ��*c���S�U��Y�w��z���@��ʅ�8u��;j�	lF��Z���q�������j#�$W2uu���|:��S��c�p=n#m��]X1�GM❣n�BΎ��_Ϗ��c��B���qub^�N�F�Ӱ،�Kn�T�� �z2���K�� S֮��ɭ�i.�ga�v��7/ XM���ݭ�M�-�v���;B'c�un{��x}tWb'���iMu��@[1�����2�Pn�Z2��>�w*�{<�z��}�X��
<�@*���t���y]<�:�裳�4�]�Gh��B�`�Gc��Ȕ��̽��#[Bt����{ߡ]�'�I٦�N�� ���Ǖ��3���p����vl=����U}y3�^��ߏ�U:p�6�����Tx�I6��EṶ�O�R�n�5]�����.�8�V�����<
,�ʌ�[�l��
�?hݙ����,�� ]�gAי���"H�Q�`)B��[ô*�>�|{��,�o�}�-ݾ=C2d� >}�!�$��Q�[q�"C��t\Fugc��v];�g�ڶ�Zvݜ�\�EB,�J��,�Ə����v�DR�n��{��̝=B�ӌ�Q�P�0[I2�MZ�������N{�L(t���,�M����\�wv6D��OEt�n7O0y�\�t��� _tutbx����k�ᄈ�YRkN���(� ��f��ɐ�����ƺ��<�s2���!��&�NL�����U��ô*���;k�,�o�}�-ݷ��phDd�[i1v��|>�;�+2��^>�sm��T����L��Y�og�-�NP���Lػv���um���{�c�{��n�<�*��}�!��I��*Y��*��A�[l]�]��UvI�U苲V�C�ݪ[��2Fz��ҩ�93��}���
�T��wv������;WV�ޞ֌p�m�	��ٻ8���+�����޵��76�.^�����F
�t�3J���*��2E<9yM����P�y��r��.e]A�S�+� _j�tԔ:Gx"A7��{��ƽ5��&�,w��'w2k��(Ĝ���ZH�,����}��>�Ƶ�o�w&k/����)�Y0�bM��o��}��l���J�J�� �����]Q4��K���n�շ�=�[�~����{�]ռk�Y�����{��xAe�[�s��s���TK�ޒz\�&6����u����M�aH4cI����|�w��ݼ;B��ӓ�׾�T}���x�wn�
D&�PH�P���͆s�T7���a���xU*��4��3&=�`�2�p����7f��ߞ�͓���6x
�.7���V��x����J�0	���EٿV��g]xE���x���ں�۳�V.��K�5,e����ۄ�6h�UX��&�������݌Bt�;�{�3�
�GA��{w����M:<���Վ��)�>�2�ծr��G(
J&� �A"��������ɦ�DJ8�m�&E���������;�+2��^>�r�d��UO��{>8�P�.]�����$F�"�ݑ<��['	ɘ��]\�c�Be��P��Y��OP�t�ruZ������}�� mn�w���[����A�R%��A�S*��\z���dΪ��UM��WwoЪ�>s��p�&J��NGŹ�y߼������ݿ
�Y��B̫z׏���mg�Am�Q�	�!����g{�ffd��n�v�+7W�w������<#��&T*86�B��U4���9��2qi~*R�Ҫ�uhوxL��]=u�6��Wbdݚ�0�.bln��u�������D����}�f#��g���Q�[BYy;WG����"�������	DU��6�P�4�Ewq�n���n{W��[b=����J���	���z�8�c9W����qx$=m�]s���f���+tto6����kp���[ �!�*��ͻ&0C���[���3��M���Р��l�q�M��r=À"���H����C�<�u���8�n�������.k�p�jz���]��01�a-��i,�{R,�nK�pk�5��������E?�.q�}�Lg��hrd����T��!�bj�z�m��!OGg9,�	��ι�7	lK��ߕ�Z����J������Ю����P�Cl�!��˳sm�^ w3��]ݸ�W��v�+�| �{�ցi�I�H7�-�N�o�b��-ޅS���󗏰��z��)U8��e�a�� ��J���B���s6w��nl�;�P͵�B�~�9{;���q�L1C%$�+���q�76߀k��v����=�;��� �r�>e8dPFXl���<�	Z!�N��vMmDܥ�w>Ѭ.$�M-���ڐ�\qSD
m����w�!����w6���/�̻��^>Óm��R�4�5R�vO��{ʵ�.B�*ˇ�$jgx�Q��VL�o+���ZT��`�����p�vh~[�8;�ca��m訅*oaS+�fT�P�
&1|��+T�A��Z��gn�V��Ԭ�[z������̘�I ��mX����p��
��\z�Ͼ dΪ��UM��+���F
�X* n.���}޵�*��>���wP����I�ޅ�V�IQ��l6�#"��sm��T�������Y��7�軫q�Ԭ�[~}�?��;��s��v�ev�� \7=�v��n������F��MtӸ��MZE��471�8��UM8y�
���{����3��]����K�b1�a*&^�oֽ�;�U� �a�}����<��f�=��Unm����D�R81�$/w6}����x�U-�C%��ӑG׎J���kc���/�s��\��1�O]Z�� k~�
�iSٱo�/�����Z..��K�x �&�$$P>x�4���~�x������aHYn"�m���ڿ �:�z1ݽ>����w�]������.^�����T�&K��!���vMދ���� w��̬q��(��oT�t[�߻���������Co&l��f�y�rj�����Q�[H����5c�n�{kn[��1�8}ޅWV�=f���¼ ���Wwog�-�L��3	��(�un;������}�'O���ͅ���}o{�(x��� �&^�oW�R�o0j����ޱw4㻩Y���ψF�)��Pów� ������r���.��^>�s|�=������@R��
�kW�Uu�uN��mG[��Jkr���*����}��pD�z�KF�fQI�g�.pgz��B�z��J����w�u�EE"���U_��t��v��%�Qn!3CWun3hUM> |{���o�}�wou���� ;_��Z�6vW��g��Z7=�[u��VNm	�� ^!�W�n�xuc)t�ә)$�fV=k��nm�S�)U7�5{�fd���.���z�D&�
0!QMY���OGE���:}�r��zݬK�Q� /d����l�%(Q� ׺���UK3��߇�{ޥfi-^�z���4�H(��6�,BLUN{=ޅ�V��Y���O�U��gtr��q��+̷	�d�Kpn�����͓�@vg��'9>^����w�]վ�w�K�X�ob1공�ٜ��%BPm��2�;TifA�D-�ҫ!'�9�u�12A5yr.�ґ�����9@p��F7�QЦ9��ɽǹu��
:WM�8'���c#�az8��A�B#�[Oiw׈��hTn��U�\oNtWjXA��#5�39��ήe��"9CGVF@]��縣�c�c"�wy�mE�.F���Yla��`��$�:���������%�ݸR���fDq���������"�]R�K/iRP^J��G`�h��{�"��rt��h�Xo�P.R����`誏��q��Kb]d��F�fۼ��`�U�sC�/�DQ�r\<�e��M6aAwU;��'h@�$����_oum�B�p9�V_N|Fj���������^p�cO#��'.�O+�	�U��=�{/9=گ`{DG�f���1�R�/K1R�̨ңL�Ӹp��M^�q�ѹ�\�3 l���ύ�� ��?Di��vx7�W~�ܥ���iDNt2y�f�M�+��l���*�Yb�n6����b�N�����;�����E�u9��%��`ي�'Rk�$�(? 3�{{��+ק�����y�|Fs��i�lyE�d�]�C�;Ow����;��ZPrS�T��H��W_oNI=�sy[��!h7��U͍�v��=X|�k�y��^���;=}CƝxF N�z�w����Ӱ��Fv{n����YB�+G�k"9�ߕ>܇����Z%eV�-�i�E��
<�E����ixL���!���ѸvM��9�8�
���Q���,�a��L��j�y�ϛ{G'Q�\]�=]�9��<�a�$�^�$�^�9���(�tb:�� u��{z��l��<c�S��=h��t�Me��i3���3�'=K����m�ɶ���c���-�����u�:c���;<r�n$���py�\;	��B��V���6ۛ�Os�7�!�U;;��L�L�v��1@Y�L�^�1���8�\�]�.l<`t$%Ӧ�$�����\�;�׷�h����=q�*�8S�F��g�".LY츂��`�g����9��W�vy���b�99�\��ge�0u�S\�;�� Gg(�+�&Z�m�ێ���eGt�lQ�9�n�ֶ��W�Yl�v�u����q��W��8N�2�=���nwq�\v�w��:۰�NӶ���mx��/�����띉s�o|����=�F�޺�����Y����	��=c͌r�&�q4u�-��;�
x܆�ɋ���[�b�qF0Ƿɞ]�n�;����N��x��7N+��E�k���|���c]�K';X�g����c�����E�tM���Z�7lCf��v�熧�;[��n����ŷ�����3�{}��>�˰���ۺ�s��m������}��c�S�wl��ہ�/`����n4C��s���iv�q0u�V�|����F�q�켎��a��Oc�K�aO�.K���-էcl��5�b�s�Y7nB�޷M�<@0j�6���r�Py6Sr{r��sDgl����[v�	�au�%ֹ�����x�8��渵����m�]X䞶�A��Jz݃N�6!-v{!lq�m��FD�gu�Kp�6UDK7d�����d`�
ݗ��PK8�O{/8�e�q����g��ڜGܹՀ��oA('/�su[��v�����o{ �{-:�9��[q��Um��v{tu�![��J6��ιa��m���:���;Mv�[ ��mŸz�Ξ5K�dJT���'j�<i�m�H��H�����d������>�Z�,�6%�"
eKO[��-�p#eF�&3)��':�|<��`�Y��ki:BĞi^����H�ۘr���:{��8 �~�黔�����h�8��lСZ�_�7�������Zڅv[eH�3��쯩���лq6i͘������--{�3��|{���3��J�ڐH-�̈́�����L`�TjR���dL�k�ɭ*vU5l"G�"����)�`�t.�`��99����ӿ
8Fnc����f��)���>��xL����<j�n�`܋����"���/gh�G��2���p`�oH1�9Ai./�w��ri]���ݳw����Zk���Z�.գK��ǌ�Nv�eC�]�,��X}�Pg��Y\B�1����A���l��*���,pX�{j�B]]���WG���WN��e:S�r��Ӳ°S2l�ܩ�L�.��"�d�~��g����8�����땘�!����s�FX��c������������p?m�8j(`8������C�No�PN�1]٩mە��P�s-��/-�A�z����L��G`���ֈ���uZf�{������k�nc�.Nk<��VI5��bE�7	
A�CQ��nf"d#��J���H'2�YI�n�}�:aL��	�
Ӗ�L�F��P�i�u�8*����U��\tm؛Lb���ZFk%�Bζ�%��3�`�)i�
>n!3;q㈙XR�n;v}FF�/��m7r�ݒ	툻��[Li헅�k�=����-�k����;7V��W3v.�x�W8._e����7%W`wd�vl�`��J;t���ͤ㮛�c#�����*����kN������5qC�L��f�1��v7�ɓ��v�g{("��:��O	�/6�B���lݳ�{L[�u`�s[�~~+�l,b��������s��e�u���3��Taヶ3��s�L��]��g��z#�SӲ�_�;6ߔ�E*��������f^L{ޥf��;<����)��Pӆ�Ż���F��s9f������ڶ�N;�9�@M���8A��L6`���q������J�׾ d�*�z1ݽ>�����vr�m��2�FI8Wu~�|%���Ij�
UK0j����o��2�w�x [�	8��e�Sj�շ�z:-ݿ���`̛ɉ��,ʶ�yz�ͷ��ÇX��т�P�f2#��z+���Fn���۱˹�ɽ��a�Ŝ����I�-�(���HF�����]ݼ;�7oa�{�W⪹��S��&d�s� �[EApZb�m���+��1v���^��&�kA��9��[�Ԉ�;�=�e���:.��,�����y#���L9u.�.w�q�{mt2�1w��\���<�>�|�4I5D�	�'�M?j��<��R��������z[��MCd���L]͸��J�ն_GE?���=�2��>���9�Q�a(�a��0�sV���:��-U7�9]ݼ;�s~�|��{ޥ���w޴��
Nؐ��,�ݜ]����w�fV5���nm�S�)U?�������÷;D�6��Y]�o^���0g%G+��k�^��]����m�ri�~����]͸��Vn���:<>7s������tZA�bE�E��{�����N�ﾬ��w���ޏ+�����߀Q�Ջ|=4"\"D"i�Ź�)��2i�M������� eE ��s�L�z ��򹍍�ŗ�Pk�XD�X�sq{-�Ok�.�aA�bz<̕Jb��7��V�����Ƞ�E��N��յ�|�.m���H���D"Q���>�L�G�e->�
t�w|��� O��'	� ��A@�
�wY{���� ��W6�k�j���fd�ѓ��F��"��a��d�\*]:��K������v�B��Yf-�-5�ѣ	��_!���V�ȧONLɫ�=U[��g����{��<�	�h5��qsm�����L�G�����X��q�Ԭ߾ ^L��K��M�E�D��oP��p�t+��&;�qsM�������d��,�{��W�����m��o`�UUMr�92V����k��S�s
���j:Ź�d�v�o>*n�%2�cs����՚�y��������у��;�g:z����}��G�8J�-p���R"�"(E��`����w|�2j����ϙ2B��H"27 ���v߾���31-��gv�ׇ�az�pD�n������ڻS�ڀ��mM�����n�K�mHk�7<�p�������/���Cn�&'}�|e�ǽ54�.�An	E&�4�Aڻo6<���2t��.��{ޥf��,o��	����4	07���������ǽ��� +[�|/��{��wv�{��M��6K[���߾ I��kU�X�uN/v��oj�����fϻ�iXE).38四o5�Wo��z<�3�z��ێsd�>�=c�>��Ƌ��>e�vf�f_��������j;�&rd���ޓ�x#��k�/kD}���G�>�Es�^��dW�j�;8��d!�V��|�����S�׸�^xN�l@vc-ż�FE^������*��k���<4����a�vk���b'v�.����%���6�\�`&��n����-��Q�.�`�S�Z[�=�g5�m���۶s�$pH&.����ܻ`�s����t=�L����m-�s�����7��hU�nG��ry�G��nw.�g���]��;G�kNo}�\����F��XƱ� E$�*��6�l�uң��S��c��;m�!l�]m�Nu������[�̇- �^N�Y���~����[���]ռ==g� ed���v�}�l�M'�P�5wV�X����ɏ{ְ�[e��T��ؾ����(��2`�L�I6�[�����o5����fUoG������]�y�ف�q���M8�no�U�����ޟz��ۇ��]������{M�ޯ!6r���R�vN|z�wg��v{�1�{Ԭ�[x�wwo����>l�@9c2��P=�Bcu'n]1��n��J�˲v^zG'!�	i6�4"@[���g~
����76�k����<�{��wv�g�/�e�� ��۷�J��u�dH��}�v����<+�n+]��<w4C|�b��3��f�l�u�f�{(t���ӗ�mf�ۋ�Y�6V��ȫ��͞ՙ��Ï	�I�H *�d�6� ��(��.U�`Z9\��J���Y�v�{�.��<�
�����p���!8M����oyׄZ�o69]߇�'ܽ�1ۏ{Ԭ�[g�R�`��l�K�6����	��`̛p��
����w�o|샾>*ለ�0��Wuo9u��o�|��Xr��R;������ݽ�������L��Q��08R\3���ꝃ̠�����v���c��'�u�+�;L2��jI��mi������u�-]��ï�+�P<�/�?hݛ|/̗!e8`��i�ڳum⑼o�|>����`���}�=�|]���/d���2D�M�CI�Ż��<��^wX��>���n���^��|~d����	�#�����ݓ�dn2.p��,-��Q�vn#���e��Y�<I�rgB���nS�����S���ux��n��"�H�`�&(�رEF�0�Qh� �~=���),X=���a�l�����T� N��2֟?Qt���w��}>�j��?yzl��pX%8i&.�GwJ�4��c�֮�;�UJ���wk���IK�0*X�ݞT�m��듭�훝=����y��On�n��j����+r뮹���}�wktr��y�c��31ǽ�Tf��t��I���H�Wy�+��.�Ͻ�wk5{�p�,[�_� N`�x�0�i��j!��f��.�GwJ�> l�R����R���= ��'4S*����=^�\:K����������e�V1��a��r�йC1�Z��	�6�ń�ejzઘ�,]�}�s����j�#�u�Du�9������(̠�~����_1&0Ѕ�Q�(̌��/��ILQ)˳&KLDb�k~ݙ���~\Q�>���e���쩟 >��b�V�������xf7�U�x�$�q��14a�F��:ۍ���u�`V�ܐ��m���jq�g��8VX&ĳ�1�.��UJ��ݨ��T�(�}�28O�6�D�ػ�p�|U߇�^N�z�.m�]^n��׾��埻��D̆b�$����ޥf��/��~}w8{�e͸{�*��蔺	Y�B
vno�3����]�ʪ�gu����}�R��m��K��E�� �I�n���w6�� ���̬z}>�sm��mݽ����FK[�䅜�f��v���ͿbGgRR^�mH��t캬&�j��M��ݥ-t�%�:������)�wM�y�0\[i�(xgsX�m�=Y�����>����]qmlSl[��L�7ď:�u�%��5�7n��m���\�8�<q�+qg�]. �mq�<��,�n�����V�Z���	v��OZ�V7gN��'d
���%x��}E].���nW]�VwO;��۳v�v������>Sr 9�p��8��݅�*�^����ts�{,T�;�6+t�M��CE��~ή�3�1�2`�HdXh�C ��Ϟ����w{�q���� ���$)�n��\�����1C�C�6��Ґ�C�(Ta����dӍݥf���;�?| �̝>�����=� �0����=������}B��z��������ی�^}W1�\�p��`��)���oT���v��X���LN��̫kW����x��p��E&Y���߀g�yfe�ޡU4�wiY���3���c�{����e4��.��<�*��}����98ީ�n��*���� ����	�	�3!C�W��5�l������f��un�q�u�-sP͊i��(�Ai����54ݩ�"�ۍ���wW0�x����?�����J�a�vnm�S����~3#���k��˞���'2y��'D��q˷�+n7��
�����t�:7yH��;6d�\�-?�����/�\�C�@� �M�قba�DW�t�wFi�LI$e�3���CW�{�Owvyw�7oa��ǫ}T+yw�z�	c�*M�$["��N��32�=�w^���T�����o���ۻq��YFM'�aU�_�����6���Vn��S�E�����;2�xz����D4���e]յ��Y���>�<���U���cٕ�  ���Q�i �On��Y�Og���S�iz��rD�C����{ ��E��$?��QMa���Ox�wo;�]ݸy�W���ç�u)w�<%z (JJ"����|�����vy}�n�������o�~9��|Z
aȀ�L]ո{�*\���	�(�B�v��4��v��6G��n�
���)!��$4#�)�~��'��ej�M�Q�7,�.D��f��<�V�u�!��3ĬZ#�_`\f1�ߗ�Kv�K|z��2�B7�w�K�u[6e���S�/K��fޜ����x���Lv����w��-܂l^��黗\�޹�9�jka�HQ�}6*�����%�M/��P�#���l{�F:m��&�i^�j�s�B�#bf�/������+���o5�_l,� ��s����y�/�ڈ���I�\D�y�s�ō�v�V�!ͩ�
�Yغ����'�egT}��������9��ck��.�����h�����&Ĵ����-w	�]ݜb�˸]qcY���{�%�.��rw��^q�f�d��	��X����ｚ�{�D�<��U�抉7V�ngW4c��R�q����Y�dd�^�Q.ukc>��{j���L�3���CǊe���`�~U.aw���vh�,䫓��ۡ����+�.��d'�c�������1��|{��'�I�����Bh���&�/ E���oI� �|F�9�K��xZl&�	�'�I���F���(��"e~۵msx0=���9�Q���>��⶿B\�#��?b�G�u���n�y*����v��\�5vvX߻�,�ץ�N�<@�d&,}��њ7vg¤�i������ѱ	s���d%)�S����k�u06'������}]0��s>�Ndv#�����Ur��L�����Ц�3��n��Q*r��3ʦ7)u,�}*'Cg�8��g�ɑ�U�� �X�K��&]P�y�v�{����6np�3s^��d����"��6ߵh�FR�D2b8q����QO<�hMs����B:�y�rO�^��&�ٞ�z	�f���$.gn��b��aٺp��qR����ăg(����,�Z���%i�Zՙ�6�����,��;�R����@�!N>�۰�n��r����I�g�那�y���o�"�0��:�&��"#���.�5��q��!���~Ǟm���5��S=Y�`'B҄AL�h"��Tjr���U��'�G:{�a��b~=���� [toq��p�ʎ4����w��ڵB���`cGdG�#^ݯ :�!,cK�b0銋9P��h�PH8İɸ�v��Z�U�4��>�8�*V堞����"��C.��1uH�,ж8�[�*�!���<�4��N��>G��/��A�6����:�e�v Gǃ�`�4b6�}�w��۹�������BN"t?[X	\�ph����T�M3i|�!�O��7���s7��M���B�.4���ۚ��/c�x's��{�$c&zs�u����4f���n��w���ɷ�Y�6�����:q;����sA�9^���
"����ګ�D`��EQ�m>�b�o����{�o*���n�4�QB�X��)Ǖ��RWݺ2�5���}/ۧ��@a�N�b��x�q�X��&�L���3Yf��	 ���B,	�Q�}�J
���\B�r�g�v�w���p�H\�P�0�AL]����w�aʶ�Ox�d�N��7wyUB���'�f�ދO��؊!-�Iٹ��mp�wo����ff?����{�q���=T��0:�q�J)�P8��Y������#��+�r��9W�ɣp�ZmZ�dZ ��n�dc�{�X��p�x����r�>�}��:�*�SݮE
\L��J���X��(V(�z��oT���v���|32|k�A���!�H��e]յ���nm�\*���]�V�Ywo�z������\���I�"�H�no�P��]�1ݽ�z.�������9�;���Ԕ���aU�3]��Qy��G,Ћ���\�oe�JNF�d밝0�&�a{�Ok�"Lmc;�r���C0�&添+g��7��7�/<tf(��TR�
l(BfE44����D��D�ID�A�D�׸�{'_p�����P��h;Wo'y+�����`̜q��+7V�)��v���o�(!�L�Xl�Rv���î71/lOb��=�yT�d��>:�.�sb��a��pT6�2���wv�.]fn�gu�}���%��U����)��M�Ce)	Q��{~�=[�!�����O��׾�E��y�U߾2w�jL(%��(I�����~j��*��> }�ǽ�2mǻԬ�[}�0BV��M�$\8�w�w����o{�]ݵ��Y�� �t�f+��em�Y�YWuoOu�t���w��+��J�z*�z��n�������+��5�hV��	e(�ή�p����!e+����l�Z��3�8��JJA.�oL����=�%6��W�-�&���bAL�ف�s8Ϡx�Pf�s�c��M{1��8��*B/-�8^#�:ٹ#�FMVt8����<�����uۏ�3s��l�uXl��%�z��[
W1�)�CGZ:l����lAÃ�]ir"�����nwkOV1k�=��I�4����n��y�k�ϳ�n3�Z�zc�v67D�Z��X8�����s�[�-�f3�kG\�:�V��}x�ǟ�������
eݸģ�!7w M6y���y��|��/G���m�����]�B9��.엷O#�V��R���03b`�p�q<�|�ڶ����]���~ᙙ<}�so�=BIE��$?��QMY���N�E���N��wm�x˻V�.]w�±��xJ�`� ��R��J����}����,\͓��|vn�:�Ta� hD��n����L�x��V֯/Y���_�w��ӵ�K3-��!y��np�&!&.��v�+7V߀�s��F<Ǿ�E��y�eݫ~�^����&c!#,2\	�\�]lzm��/��{?a��L��h����k[,����X'�����o���v�owv��X� �g,��ǫsd]�&�MH�(�Qgf�ή��>�2%x��d�۲��o3՗R�k!WE���U^�fP\Yx*M��W.���*�����w��U��<��P{�Ϗ~?_��&%�D���Y`#�����y�ִ��^^�sm�~� ����(�M�!��P�Y�o�ޱw6㷩Y����3��fd�s�wvy}����eC!nF�-����/_����{���ZY�UW��>]�-����q	�J,$�-�[j�B��+��}]v�o���r�76߾����@�&Q��l�Q�"*6Y,J�u=u�����B�F���w;�.�؊u͗7k��,g��x���Wwo�u����Jχ�f�]��O�&���ۅ��0G!p�dgv���2��>�^^˛S��.��y�k�@n��;�e'P��bBR�n�9g���7V�)��[�w<r���
n��	HA���W��d���P��GF��r=9��@���E�VC̃:��G���'9U���zz���;�;J��&;T
�(}�m4&��(���|����軻o��.�[��RaA,4�A0�M;77���Wx]�K{�URӻB�p GoR9k��Je�IA�F[js7��@no��<�V扞c��Ɉ&Ho8�:G��dN�w=�c�#jN�q����b!����ֆF�(�����_���jU������>���7�f�i�.����� 7������UU.;�^ M�(��0Y��2�j�RZ���w��&|>�vw��e���u��ބIሥ)#c^�	�|���y{2�͕F�G���k|cԊ:*᱄��]`8�u]]*���V�T��<���z�D��B�7�������PӮ�z���v���_M����T�DR ��RDRF�|�ŧqy�]Q�0���a74�7�ݛ�|>z�瑓y6��3$��OwvtW�P��bj6��Bz��'X�ܾG�:ƪ:�b<�!li67�!ח��=r�Y	��62��Lf<q��+7V�K�����}�ݵ���v��p�W�Q-����Ͷw�W��M��owv�}B�Ӎͥf� /&N��^n-���p�qn���wv�owk�}��z�윛l��u����YP�$�m�a����}�>�?`�t�7�Y���_�E��| �W����z���BlAM�l��GW�R�/}��}���1��wv��
�O<��^uS{(Ә3��|Q�v������f�M�V���O2d:nNsf	��Z�:r.D�.��;õ	�N���E�NT�����i�t�m[����]�v�AXB��`,�Ð2����)8�v*��u8�<�v:ui��ܛO�[�zSD)nSN�q�>cw<n���n4iF��1�Bٺ8��DnWj}�m��u.ռm�<ɧj<�&z��sۊ�<���l��P���퓻]q���u�v�.�;d�F��.��^���u�Eэ�Gl [�Ev�V���p�Ρ�7��۷�{u��\�W.]ݫ���tm������O�nv)��W67n+���\�/k8s�t�(��D�r�[f��i�[e4�mQ�[}/��[�y��wv���_� f^J��\��z�H��P�0����y�U��fO��U:q�Ԭ�[y3˧}T/����Z��A�9�3#;������ku�χ�dή��wm�A��w;�`��i�0��۾�'�ְ�[{/��n��u�������Y�o{Ԥ��H4�A0�I���y��ڻ~ 	�wv��
�N3=J�շ��9��+I���k�.vt�w/G�n���S{8e�7]���j��d��H]�r�-��_�}�wnowV�-���ɝ��v������ш�
4�v�s��7_����s�|d��Og\`��ˁUA�'s^}�a�����)�l�cZ���o-��u^s�fx��U���)\9F�=*�E�]u��;9
�赻*�~v�V�U�Ir��˛�)&���o���[�y�b���fd�xF	��!�i�ʻ�kWz����|.׀�fL����z��۷�$��n`#���u~3���wo}�wnoS���>�xy{'{� ��*QF(;Wm艙�� �{�1��R�um⾞���¨w��Yi�n0���z���g�i.�s��TԊ���v8��b6d�L��j	�c2����Wuo�\\�y����<�|"feü*5�BÆ�Sn�v�����^L�@�T���ۇ���|�ޢS�E6�bB`1���y�]���D̦k�g?:�s��e�=rgx�v�ET<�n�qB���s��-#��.:Ä�5�f�E芳4���A�U�����Mnv(�L�_a�;���r�(�6sN�%p�$�`��WH�v�{Ԭ�[g6�sp��rSi��w�*���9�l3��{���\\߀g��ڪ{��&��� �m3 ����]wmx�{޵�0�O�5U=�����T��P�ai�\i����)[Q�U���X\�sûV�B\�)��b��M&�̬z{�.���©M7x5{���̝��ݻ|}1�[D��h��-�f���'�|=7;�`��7���g6��dίZ>���0��V���Wwo9uݿ}��=�ZÖ�����9���d#��1A��ڠ-_��*ޞ�\\�gxU:�Ό7�]U4zUw7f���T�����O<ZN��`�9��̍������%�GB��jihSxW^Ga�D�P(=H�e����-��m˜�뤻�ҒDM|���6z��S�I!�A�4�ݸ��Vn����^�j��u��������P��=�i��i��Q�"���D������ [j�8��un��TG�z^y�m�[	4J��d&I���l��S�n�j����������{��nl�w�[/bJ"���j��u���̘�w���z{�qs�s�ў �Ͻ�ޘ���
4��������wt�9^ ��^�j��p�w�9ʈ��
6�{���W>���ɶ���ڻo4r��}��|�wYÃpa@�-(Hh�ӎ�����;���T>������ٗ�Wز�_��I ?8@UUK�j� �I�����ъ��}DI���$�$ IL$�I��$�E��A`B_��c_�	BI�� ��_����g��w�(�����h��o�����������������Q�߲H I$������O�?hI&��I?�'���|f��O��?��ܐ �H������穃������_����HO�H�d��mMjm�m�ږ�M�-Tڦ�-R�M�5�mMjm�Z�jj�Zm�mMRږ͵+fښ�mKi���m��fږ��jj����͵5��6��6��+SmM�U��6�֦ڛY��l�R�Z�jm���mM��jjٶ��i���fڛZ�j[jj�Z�T�SmKj�i�Mjj��5fږ�ڦ�ղ�mj��5�R�6���R��+*�M�6ճmM���M�e��i����jV�mJ�m��fږ��R��ԫKl��jVʴ�M�5SmKjm�j͵-��R�M�m�5�m��S[l�SUSmM��mMkM�6�MT�ٶ�֦ڕT�M�M�6�+6��Mkfښ�͵-T�SZ�l�Kl��ښ��R�6ԭfښ�m���mM��jmT�M��ڕm6����*��R�fږ��jj�6Ԫ��Sm��jV��ڕU�T�U�R��MT���mMZ����iV��M�+m6Զ��Skfښ�6ԭ�mJ�m�m�ښ��R���V�ҫ6m��+Y�Km%m���իMT���mKZ��Smm�jZ�6Ե�-�j�����mM��jm��V�jZʴ�6�՛jkfږ�ڕ�ڕ�Y��R����mMfږ͵+6Ԭ��Jٴ�J�i�jm6��m��m�l�R��j�jk6��m�l�R��-�mKZm���ڛ[M�6�*�USmM��mK[M�6�6��M�-M�6m�SmJm�R�6�jY���ڛM�3mJU�͵&�SmLڤ�SM�&ڔ�Q���je�&ښm��jfڙV��3mE�Kj-�&֙mh�EZ�j�6�m�5i��j�ڶJ�h�i-hڴ�����oۚ��[����Գ[Rm�6ԛjM�&ڔ�Q��V��jm�i�mMSj�͵s�S��������H I$O�����F�?��7 I$��}���?�������?I�W�L~�� I$��'�����<i?|� I$�@I'��Md� �I��d�$�"}�ߴ���,��h�_�����E $�~��O���0 �K?B~G��?KT{�M'���| �I��{� $�~�?�����~��}E��1���pپ��; I$���xL����G��~3�|?  �O�S��� �O�����o�����������W��������/��#�e5���`�U���?�������  H� ���@            P       o>PIU)QU( �IJ$UT��R�A*��@���x@$�$�  ��B��(��
P*�R���)UQI'� ��n�E��GA�zho(�
=����n������G�UR�EN�=�>��eG�^��U���l;7�;���yU���u�Y9����:�ET��B�Rܠ	ԯ���{��n��^��݁�:���-g��/}ϯ��k݀��#G� �$)@�����u�����a�tdeKGv��M�
R�a�E%(��(]�_n��hh{�th�]�x�{�&��}�|:x�>�����*���R���>�`��>��|{ �9�9����w�}������ ����$����J��J�H��^�
r�{�4z}�{ �W��y&��'9�!Z�""���tgj�G��y# �d�c�\q݁��@փꔨ�y�AQ�$� 5����2u��6�y���2h4�������{>H��)TR�����=t^ླྀ(ѧ��u���dt�z��1�   ��JU2�ɦCF��22  "��	)J����d4��� �FF������UP
��0Ld�  ɀ��%*)P 2h      ��D���CML�4dh1H�@*���&��4�ɵ�h��6P2d�G�?����x�����~a$$���HB�II |�?���� ���?�������/��ޢj�^vڶ�K������@@tbYi&4���h�>?����O� � �����}ۃ��c_��f�?��O���_�J.�ػ�jE�u_�2�-�.��95^�^����ѻ9S�y�L��Y�Q��1��R��]�9rj/)�8wF�� ���{���_����Σ *���*��ȅ�HO4^��6<�dp}]8�vTn�/���Eť��JỊ��g.�sr��T�#I�+7�;�ś��Ϊ�TѷeH>'�`yAS�܌E��<U�0r�1�~K����L��p�ܞ���;\�il�7 ����v�f��x���܊r�?Qz��:<��D �И�҃����f��֞GF׽5��59m��[�V�oi�aM�Ob���!�-�pZ�|�	?DV]wG���+��)G-���C�ʔ:K�X:�K�v�	t��ɉ�"HP��&�;�X���r�	SoRw�*�t]���C]iQ���Q��t̏�Fh8zf��P6��F����'���E�޵�%6���u�Wb�4 .��k���2�/��
���9���!Z���N����GL�Q��D�I�y#�m��m�� 4�]�l -��d�Q�%�Qs6�	]ɧi)*������~��m��f��"���Y�G����!ŏ���.�ɹ@��}�j�{���ԬǕݏ�k⦽��[a�\�C�tn&�R-"N
i[�7�nS2��J]��2�M�Tx�.3�axAOj�lCU�Lu�'N�F�
�]��[�.�Yv9�d5q3�u�i譡�׺�u�K9�A(��Av	E{����`���Xn���vnW�=ݢ���Ó��<��i����������^�u�=w �n���P3��=���&k�|�#�m��.���o5�^��J�� R�T�e�@�wS�tS<=��oO�/��z��-�hl]��2m�Y<\M{��ФZ����0!>39����T��T��k5�+5��KN�Ю�ڻ��B����p�cӚb�EJ����_f󴜃����0i�;z�ߪ��0Wu�O,o�1.���s�΍x�� q�`�.��LQ���z�V�7Q,5ܚ؟٣��"���e����{o,�&N������B3����\�s{;t�����Ȝ�]�t�x� �}��7�,�t���U���jF~U��C�z%����on2�`}��	�)s(x�r�:���Ȃ���k�Q�:�ў�c��bҲb�q�W�*:0(��9���<V\�=��[��h���d3�N;�6ޡn^T�nц2�]�c*J�xs=\Оh�T-�5O�����%#�s�����pM�z�m|��m#��`t��Y�IΏfv�O�t���i����ތ�@R����On��a�6��˺U-Z:ˌxi]�gx����s�#7s��:����WVl���ќ/w��|l�c�V ��T��o�]�:Lг��7m/�����x6�2��yk�%NL,�<a�q��.�7O*�@>V��Dzw;Vnr+Bk�.�n�q���C�x �+疇�m�<*ku��l[ϱk2����m�;�<-I6cpVsl:&�|�����D�z���4=p��X��f��z�x���b�����^�HqP��5b0j�մv��vn��8̹S(#N�Tׇ)��ǧWE"@�-�`��I��݌i۲uTn�p�X��f��vI	�C�ܷ�ufMTWٽlWGL���ԛJ��9��w����>�>���WQ��_^�B�	�E�]����{ Ot�<���v&݉m�1��s����0R�E�h��Q�qi>��o[�x��s��7��KYz���TL�,x�3��1vL��^��&�j$4��+��wj�h����E��u����l]�jh>E�;rk(ŝ���R�<z����O=�Ǥ��U�:�x���s��� ���� ���}��v	w�!5�I(-�(t�z�4f���a6-*���o���ۺ�;��d�jԎ���Іp�߻7��z-�^]�$f(��`�0�ߍ��x˝�)�vU��՜�sN;��^ǵ��h�qn1D��l���Kz%��7�hc^�:\�D�T��F�+ZR����񺶗D{8쬾�'ܻRE�����=9z7�>���bs��GE6�����[��b�5vnGz���"�U˻�Z�1=�E�@�0���5ċ�5%7��@�[�)`iEv���z2NV\7��t�{v&]�	Lp�Z�%�kwb�x3��ƫ`�ow�dtg5DBj\v�݃�������ck�ۏ- ���؊#E�ټ�!�;F����m�Ǧ��I".cCF���УL#���n�ж�ABC�L��B�d�1ɪv��Y��Pe��nVK�2L�kY�.f�v�E�Ji4���:ېC8{�)����>���c��'VAē�u]����q_�Yk�����V1���LqJ�^�3�	�L\L��-X��A�_V���I�4�ݛJ�������;t��\J�E��d�yl���Oo%�o��<C{��j���<���v�JBO�À-�f�1�9�����P��&��e����������U�ix����v�ժKH�(x����Q����6A��PBk��i٩)��S�pX�;������{ó��䱞g��S�7�9�}�+���[��5�������c�h@� �7/gQx�XoY{z9�F[G�no� Q�]Z){D�`St9ˎ�,�8�0�%_)x˻�^�%�I�-zx�p�L��-�zd��i#.Ν���9�n�y�c\����N�3Km�nTu��m[WA=w�q�:�9{:R2-Y׋�����r͌��s��u
��A\6� r�r*5߻vr���J�ϴ��r���%��r���f��u`�庛;�������ֻv��.�����>9Eº��c6��"F��m�6z5���E�C�q�R���e����Wٺ�H�-u��쏏f=��NR�������~Ӽ�ٰG�#�be�:`{�E�`4�xVb t�=�}i������Z��cxpi���3Vĕ�f
�:5�
��O�*lf�_oB"�:��w`yIyy���S�c�&<�*P��rȶq!���� j:�!k�o���k�#�qkzr�.��0���vf��t9�)4����b�Xʊۆ �9m��Q3!��i�&]ǃ;o�Vs��I:�{�������N���Ƚۓ�p���[x���crH�B��x�
��[����ѣ�f�f��x��,�m�*�jdokz��0k/�=�{#�QZ뵝�Þ!E]xi���>#_u��t9�k�W[I����wJ�B�Gxu,�bk�{��ӕ *�QTCa{c��'�I�sd��t�G�
:.��Y�9V�sU2��`9e������qY�X#�7-������twB��u덞ܧ�+Ƚ�@=;��7R�Y�ELl��&��̺Wov�{	C����p%m�7M�h��v/�G+b<7��%���w�@���"��B+�b��h{f�޴o̕�ON�t��ӹׄ��&���5��SwN���]e9*�WZc�� {�|{���0Cy�ᇗomȒ�1�����ܑ�'^�;UT��j���kV�٭7 ѹ�s�g��=�wylZ�����"ǜ��M��b��ȋ�`L�v=ǔ.��ҭ�$�}��]��l3-���@���w&�C�D�b-ҭ�����m����9����O�I�t��=�Ɂ{��y�ŧ`������	���tba
(祋���� ��ɇG���mU}G��?��`���|~crϜ��'�\�����C'F��b[�6,u��;�ڎu��r�sb6�]��t�Rb7�l����D�hv#3�3c�?��)��N�j���v��m/7�.�D%�%6�[�Yf�A�6掷�f� ��i����+�Sk,�ǽ햞�Pq�d��t9�9�P��\-�e6�Ļ+�ۭqe���Rɕ�T)�[3Gm�xM��N���{]6t�_���m�M���-.9"������3��hkXG�E�ux�Q�#�,�v��;��R�g�����O6�}�(�m��fƚ�vz�(��{.[�MΙs]�-�0�(��R�7���.%�@v�z�y�"ck:Ώ\[]�m�Nq��W ��Űi�f�!����7CH����p�[�U�knm\�n8��u�{]s0���t�]�CWT�E�V�iq��Uڌ^z�F��,�ݴm^k+b�q��6�닍��3�¾u�W�O�$k�,J�[��H��,��Ζ��bV�U���f� jGT��ZTUGbV��*q������0�u���<t�u�eᆬ���K�]�t�l���2�Xn�D�*:R�,(�\�WF�6�8m��d�����n��z�Q֕8&-�$�D�	kM�铉�����_+G�/c`�mu]�*�iky��l61�sۈ��[ ��8,��:�\��v�lu������� ��4��XUՖ�Χ
��[n�4��s�\�X�ON�pX˻M&�ѻ�=�_,u�6g�����bM�[���y眉�MםU�N��6�t髬�pm����c� �+��sf!�#KC��l��LԖW]�5�B\Ǫ��BgCP�%��]���k��w�$S?
q��ghuv�|�Pn>:�&g�1V����*�-P�jD+��ƲԴ��B-^;�tՈ�+t��f-�ۭȰڶ�7Fu��]/��#Y��,��R5J�e�i�ѥk�5�m�(63%��<�u����sǷk/c�n�X��Z�;'D��ܖ37��8�[	K����=m�\�G=lI������bW(S:��+F�0��-�a2!� ���N�m���ۈ��)MU�:��Xm,:�Pv���k��%�C�ۓ���q��m;�][�d�փKY��턶�"�94%�4�F��j5��\����^X��Y�݌v�S�,�k�׀�1m{H�G7/�<ۃhzoBձ�9D����nl�{2b-[�[��eȑ ζR�l�X٨4�j �6�v��b����,�����T��-�콲�k\}�F�a��-k-po-���Kokpd�M.(��v)/���{���ͤ+��9��z�e˗Q��g*m��Ѓ�+��.���E���B�f0Z+(:�V��&m���(Ŧ1�l=��:�'0�c9uj����tt��!n,���0��Ir������߯z]=���+��_1CB�ZA��+�j�s1��=��5�}H��BE���#�r[�A-���%B64t�v��JS�ɗ�1P��sfs)e�K*՚��ܩD]e�"WM�X�� Z�Xa*�
�l�_���y#�&��c34�m�\�R�3�V�����ò�	�8��mrQ�:Xܦ������L�-q��5�����mٝsGc9�&z��y(�`�n�-����-Jѵ%�v#���'ƮK۞77��L��P�6�X�҉bj�+����	�cGPͭ�6U�VC�A��Y]��MO.
�Ϣ���GNp��pLmT��%��ڬn���H�b���3u�\5��ϋ�M�ָ�:շ+��J�^�n=l�،v7�O1>����{X�U;��1��ر���K2n8�Y�Y��ьe\���jf�r��C[�e�zU��a�O������pF����J����+�YhY�܉�����t�[
]W	���rN뎇���s���ۛ��"���];[���� *|��=�`����S��Q�� �5�6e���+�4nt��r1���97%vܜ�]��(�e���hf���fһ9,�ϼ��4�&��{g�n��L[�nfi���m���� �qe^��JF�ڱ�%��X��B6�KvG�Vh�F�X�Q\A#L��#DRj�ǫZ�h	ر0Z�c.��h�ak)*��I��K�۫T� ؼ@�� �Y^q�E�m�]`"�}��w;����v��<hh��IGk�ɮGCðU���O�ds�ݪ>����b�$n&���#�E�1K.atWK�u��[�n���J��)��ձ�R�[w[u
�7<���=[[�5ly�%�4j��n0r��y|j�%i�W����e������=�m�])_XKwϧɺ�y`;+��a�<j㌆O���7۵3�<��o�a�=��))�����c������݀��p�{uɵ��}iOj��V�xxɲw{�{�+kgOcE���v�x��͖��G:�n�3�,�n����5ˢ���ˌ�m��>^ѷ�lu��ư����%��28�ͦi��G+y�:��%h�c��,@�*d��j���뮍=^�"u�քH4���k�Kf�o
f��e`7G�t�X�֖�b����s=�Cn'������8�dɺ�rnw�wO���^���v�.��kjx�ָ��]��\u�.)��X�E�ȯ����q�0�v�r��cX��nf��%m\�eM����p��wuM�=u��E��״si��.��c<��6TW��,�K��S��<���w`3t����=t��[�5X��p�=;����Cn%b��͋��7fظ�w|;����M�է�����^����kC�����Lw������{����]� '͛/��Z���>oo�g�q��"J�5�32ktfVX58��%�N�U�
�x6�9g�,ʍ�
��D��B�r!�2�5@Ü�a錑J�<�
�l��47VX���J�v���d����xn�_;����<��l��'$P>ڏPt��{U��Q/�Ӝ�1GԹ�b����N/`�&���Hc��t�/M6d�.�������M/�:^�m���kع6C�eC�sq-��F<���9��9�}�y���Kr�D�flgnE��LB�4n����Ww���+d{�5���:�˷H�5�:q!��_o�[��:��J����n����YM���c4�N��ЮŌ�,�V�w^ی����K~lM�9oہz����/�|^�]Ow����f��>^�xpu8wS�xb'�ŏ���}"YoΜCr�Tu���g�Z�����;��F��o����Z�>@w]{�l��q�%�����y���)w7oM����=�ޣ̞�䳻�S 	��Z�q�jOt�Z<zv�U4 ׬ѽ���I���+m�ܜ��[�Ԛ�8��ݝrD^[�]R�^-��t&u*�k.i�T�\h/d��>�2{�m~8�� �����{��=��p�ldۗݔ·0�E_�θ1;�*t�sM�`e����B�p�?:g�=�9*+~䙭���yOmK%ӄTk�Sqip����սL&����l��`�k�A��c]�����{�D������UBtCJn����z1/�A ����is�k�og2b��D�w�f��+)µ�ZETD#r�eeU�H�	m�נ2_��Cj��q/Wr��&���瞄F��<]U$��j��}�.�1V��^6
���{/�w���u�k���Ǚܺi^�t���=�A���H�v`��;�˻�x�{R���w�7{!�� -���<�����\�m�t�n�9;�}��ކ{ڒ%�o���ygmݾ�j��b���2�j�z�+d<ZAy��J/b�F#+��^�(����9g�y,��`���,B�睞u�o��.^)�<f��Y�]09�1�F�.��	H;��!³bV&�dh�m��r�5b�NոU��(b���*#�(�����g�]��Y����<��h��=�>��������;��-^55۴�-q����8#1"R:����� ��&5ⴳ[gy�^�u�'���AQE.����X�s�yl����4'N��>�1�8wt��z�E�1�Τz������V��O�w��K}^�d�{_z!uCw�}���:g���N���6-e��K�DV���� ;}�N��η�.���?Fn{g��{}��>0_=׵z����+��r)�y�q�l��������Uo��С��`�zbDe]�y ��M��h��h�;Mԡ�xQ��UI�CnF\(�ݍ{۞Sڽ�.�|��{MΝe�����G9�l�=�����Ku�/ps��R2[���M;����k��J�+�\W�ۀk��>�nL��ǸXv���g��ǯ�4���c��-̻"�g7{����}w��[�=�G7�n@y�_-V�}3�J���9;In״�⣘rv��TY�ݟ6�%f@��=�uJ8���Ӆ�d,���zu����:.�I���eZ�Դ֚vS��;E�do�28S0dCw\��<{G����f-�S��[��Yhd�I�&�`y�^Z3��������c>o8Z/��*�_�Uyz���x��=�"���=9j���Qҏ-bֆ����g�m�t�������,����q��9���^����l�H������d�Q+n��;:���$�>���n�_�J��7q�H�7�U��iP�K^�=��1��:�;�r����������S5~��� ^�;�V�/oe<C��DC�Ta�٭fܽ#sl lA;�˱a�����ې�U��}��'��U�}���W��������}�5Fa�{�N��	�{{��������o���/^����S�u�{��^>���bN��N�-���z���#5��%�I�O���Lޢh�ֽO�^ὬM$]�.�U�xl��wnǔ�<@�:�NNIf�X��J�V
y}��~��JT�g�]����������E�s{��w0=�/i�dI��b�*^�����[�;��ΣV�'��kἙ����G��`������>'{�� dzw���\��K&�V����*pY��3#Z�W�^���c�<<Cֻ��z��s͞�}�_eǹK���+�d6���n��dR��[U��3r����d̝�q���}<ג�]�� �$��Y*#s�Uݾ�6\�9�n�|�
K��*-�M;2Ė�� P�{��բ�)��jQ��Â���qۋ��5�v�Y c{�xog�^QK�l�n���yaȰ4^�S
{��`�u>;�8��
�30\�V�NP��)i3q��7�FNu����+�D����v)��D�̒�#66�kƚ�<9̹3tE$���N�i�t�M3W۾滻�nz�^�s[�7t��>^W	<ɷ�C����wJӋ��+ch�S�W$S8������f��mC�M�b��2�S0n�S�P^�y[���6=�tX�ɐ�	fw��ϫ�Sğ�}݇x�y���Z�=�Ճ�.Ժ�����������z	;�6�U�c}SF(����c����#�m�p��q��#�8/Lh��������g{�W�=�o��ؽ�����47w˅����>�G��j����v�pL��C^^]�����U7�"4����OM��T|EKwl߆j8}'���!յ�{v	��{����՞�����ٰ�`�'���&�ׅ�~7®�%׊B�������['�e�o��nj��v�w��@t-����U��j`ZN7���M{�BR5�i����%����#�1��|�()�7UkNf�]em�e,���vO>��d~^��=�{�h����wv5�+�ި�o �cbr,$�l�>�XZ�+��>��Y�oV�X�w���fd{ {x�܍�P�`8�D�ӃN��t��>�w��#����ŝ#E՜�%��>^��y��=�����ǣ.v︲��x��z�v�0<��z���t���W��T��S�ݏl�����S;�K�������w�ztc�+�L���{�/��5OZ�r�BM39�����DF�جZ� pXD�;� /ČDf����L>/���R9�l���]|#�+���}��ƇY���k:o���}[��
��ش���]�/�[>(��oE��E����\�aX5�yKZ���L�W�%��z��i��c��G�T��-�xtf*TޚR�LE�B�dFQ�b��bꟻd�����ń�z���\�͚�ļ�;���>�5�(NN
��ֱ$����U��B66��o����f��x�B\���Yץ}.��Sú>�Pz���8Eg����Gce�@aݠP�&wV�TyId���`#/	ِm��Ĺ�o<k�����nol�8�)�i��vN��l>��.�a%O=������5��_"�mj0�m����؈h �ǪoR��OA�5��x����X�T���˱��D����n6��!��y-��OMXS�Ϟ� �����"6��ݼ2�mՊ������q�������ш�w��������Bk*cA)�}���w�=������{�7�/>������8���6-a��E�A�T� �p����LO^����������/��م�
�}�A�+s�����<�=�Y�sF�c�^ BH����#i+Ko�Ͻ��ͪ�c��%|����b]//g�9���+v鋞��s�f8`�N=��C�\0���]#�\��g�g;s��#��V��`ӝ��e:�q�Tc�J�P���H�Ϡcdsf�E�m�e�l����-Tt�Ҍk�Aq�:�f��Dm<��Վ�l]��S��</.���c��u�ڕB�c��÷���.��;��=!���b��U��[-��ݒ��A.7lu���Ū��6�RSJs��V�PtT��E����^�ŮC�>�ݤ�ԑ�N�6�K^d��0Wp�����TL,v�-�t�q���X�8��k��m�\�Vg���b�f��Pk��g>�s�p�g�:���S��-�}s��ڭ������Ed�5ٻF�١j��RiSd��^ΤC5�Y����lb��8j{f�6dvy���ѹ7csQ�GW�N�\�2��.ÓL��T�j�9�j���r�c0e��J`��M�yM���us�ג��Z۶S���cp�Aۛ�נ� B���(,��t�ńV��`��QE��\�	�qA��[��R�v��md�ugn�\�Cf��6��1���~�D��$��MW�2�USM�sf�(��i��ɛSq"��!�Q��'6o-2F�#xxe���>^�  ��x�aӄXſ �q1!ZFS�B���������;��J��d�Q��{�,6D�+k�9j Hw4�F#��4����#��NM ��z �v��G
Z���r� ��l��C��fh'�d{�b��_CY���^n<��'#�	f���MW�Sd�ä����(�jF�J:����^p:�b/�y�&GEE1�bF.H���Ty�)���	�tm��ySV!`핗���;�v<8�C���O� �Qxu:$85A�� �Ӹ���Sz�&��i�������\�y�n��j���H3����	(�片�pkb� ��C��b�}s�!���2s��1i�E�q����F!����!sf0��|u�O{�h�wn��6�F�Z2�[�ۍ�{e�ۈŰ�"l�{ֲ�ʐ�qm�Z�h:���zoT�+�-��#�(hm4u�)Mȅ\Onk�.M���谚fX˳.ְs�Es{j�sx��]^��Rn�]Żm{u�L����۲�3�I�����^E���'>����C�`6#F�(�h=h-����oID���3��������4���]�̼��aQW�%q��e��S�cȼ�>�&cuc2o��S�Qs�J.ʌ�n�<oWF���P[r�1��=��v[tM�d��G��h��رq�´uVgm�&����j٨���ytE_x
�gqw�R��i�=�K��$ׂ(�RE�Ě�o��L��Z�L��ث��;kt�[�==T����P��U<�㙝����ـPlOF�Yb��x֣��ރ��\D����!�e��,���J����2f;R� ]ܹ�c,�����D<�Κ�9�nڝ@d6ѹ��n)��m�f��*��C}0$-Ģ71B��(�Sz�3�TO[qZ�����%5�+���U�=�xn�!zV��2�q�k�xL]��Hu�;M2ˊ�<�M c�qP*=�C�������ﯮ�s�/^\���.1����-�%fm[i�(�9��{����V�xK	�����
�����f���*�q���� ��	�Rh�Pܼ�0�b��GJ
JG +�y�&:��z��wO.q���i]�9r���V��>��N�L��;���y��j7
��="��EN{�5��x�RWBЁ�&ƾp��3�{#r�U�r�
�؋�\j��h�"��8!���Fp\K�㎾z��en��p�.o9����.*���Ag�4���7�!��t�Y��5�Z�%-D�&[D��v%iGUo�&o����e$Sfb��&��^����E#%����{���Y��&�,9܏r]�l������l8�����zrحűV�(���r:!R�����V��Q���*c�&q�:��HYnv6z���K�=��g*n�ǕǾ���"Q�T�h�F�msuu�*��G�k)g�5�qp\v�v��I*p��V��JA���.lŀ�j���:l��Q���ۭ8��H��c:������i�9ڳk��gus�@]�sC�?O� <x<q�N(C���-�e�_x��V�J��ׇ֞����^\��;6�L��v�T�f���ы��
M$���b�aTl�j�E)�JA�}R�sa���I���PG|���ƮUG]�����,mANLWcq���H���ҍ����T@nh��7Z�=�����.+�*�HC�N�n�t���E�7Ѻ��%�"Gf�{�J�y%����:_^��f4��s$S���=��P��gb�9�;�ߟ?}޼ys�D7I�D�D�DiE�g���#����R㸡��ބ����A8�2�����j2�԰x���H�ᴑJM�@�r�ҍ��<GȂ�ii��cB����U�Z�9��YNE�jQVC��{&�9}��-��;�Ff(��1`U]P�H������m�uV����L`�ڷp��R��7c�Kw�Э����39������(��$���QkT�Q3�RQ%�ӝ�we�j1\V=r��lI��Fk\<6�h�X�����w������uî��ӝ�f�&���Q�F�Z���c���7��t�N����x�����3����ݶ4��*��{�	���I�^��*��xu��DmR��6RP� �j1VT\�L�dx��i��HX�
�R�Ұ_uݢ��są']�s9'��,��L$���L� 3�0`�I%4��M��t�=�wr��Wx�z�#���J�F�EC&!�\BP1@�7=K�C�j.]�Ü2����n']|=����]�jq	q
c�{ޙ��b��}NǤ���B�����k*�� =�Gf7:o�Q�T�x����u��������h��#�]�[�+J�X�e��[�k6�zt��C��S�MirG�ngjT$��Cp������:vK܌�5,r���k�WU��-��z6�nի�Q1�Ks�L^v���j�؎T�cK>��ك����[<=�.i�wY�Ԗ���)���6;�Y����¸���]F�� pw�;���q�ِfhoNE&�p���?'��@�Û7�va�u��f���:�u�k�0�H����[YV�ޒ7R��ؓ-�Qsq�G��*'����9�}��-�]��f-��cw����2�)D��7�.7]m`���f.�J(Ia����rN��rSӧ|ď)�w�K���v���ilokQt����M�i8h&Ѽ�U��w��f-��u��q	�a�V��Mɐ�v�xIs���Gi]��,�v֝��QH�)��}��뫧��2��b�d�&u���߮�����wϟt�L��w%B�x	��b���!�YI9���ȼk�,�q��јQa4RJn5��n>��q�ގ���X�	��SJhܷJ�`�q�ً���&�;|�_�v/��ߟ��{j�J�7�[����Y�|"=&��x�RY�%#��"�L�s��YQ?�J�1�0+�7�VF���`�fir�VϽ�C��L7�mw�}�)��{��¢���L-{h�&�7��w��Cbr��?nr�Hy�g�
&!G_gr I�n�֢k'���TԬ"���^��mM_�����F> ��=3��.�U��if�5�ՕNg.���9]Vf�@{�ʹp��q1vN���ԐɡiG^,=���]�';���-��)Q�����+��,�	Ngl�Fx���������\w�8o?H�����B�~Ҡ��=4+&n�<2[��i�y�Q�<�uws�� �o:me�݃�s>�]�vh�v���DJT�h���E��J���V��-�ؐ�T�e�,h�jwp�Ț�5ˍ��&���}�]4DL@��2�G�v��(��.���!����0"�^L��p��ץ��G�?W��`�D���1h�L����gvPc���<j� g#�2"�;V��
�9����C(�I�Z�)m�&ݸ��%�����
,�.��Tp�� N�mV<� ��<�����G���%� 3��XJ٬3�(y��n�X���NY�00����E �r�15�[�S8��%�������.h�3�6sr����d��ō�W�F.�VX���#&���Dc�Ł �GwWjX~	aH,!4X�)v���>9ad:;�c��ӓ9�;�,!�sơIb3鲎�i���|��PK���l� [7pG��Ų`߸�7H��n
�Pl�dH�	H��ō�j=�e�$-��.�nU���T�>B���#�sWU�f	���9����R��)~������S�y�Y�f٪zo��f=�<N��m���Q���� 79\ӯ���dOSq��Cj���=��v%Z��o�nӸޅ���S�c���r��ݿO��~{���_}�I֗^���R�(Xi��n#�S�N��M��q�ȣuM�r�=� �l���"����\<8�;�_��v*�x@������2�E5��E��=^�S�ӎ�EW�2�%�+}��f��Q��kjb�*f��\��ܚ�M�D�3N��������g7�c�Cy�Q6b�6���	E�l�F+�xޟGwuv�������K��+��jI���鈸.!DQ,�D�+�#!�oFke����v�����,6���sy"c�x�����U��tHc�|�H�H�w�~��k����B�uλ�IS/�}t�X�KH��l��֣��m�)�����P�vf����ۉ�w{uK�Ww0��/��	jͥ�%iE���>��4^<��%ƭ�R��wƘ�֪�8�uML��ا}M�p'W]f��RE�Cpp�)�p�b�"Zi��ב��4e��\ˬ��^l����밽BU�<���v<�٭�����랂8��샸�n�95�u�ls��ZC�ƃ���f)�&d��\��ilj»��W�ؔliF��m#`��LciLb��.�S
K�j����&�˗�:H��)5	��_fPa}/����R�AWĝ��)�e)_Z]������1�ҷ��+��s�\uV���wg@�/g|μD���������¾ާ���c�+�0�/>�c�s���%�1�K��	��}�G�M瀽Y�i%���M�3&3K�1�j�Gkc���Ϸ�"ZF��B�t�W���{�3њ�}���Fc�U�#����ގ���e����[SKO�O��M�lK���1�Fr���߿>os�=�(��B%0�14��q�6��l�Jc�2{Um�T_P�${[�dw	.\ww�oU�W�{��J�K�R�Re�$�}�=�tdƔ��s3�<<�0�bϒe�Kl���{��ٖ~��z��}�Ј����*�P�m$뮌n��ml�+ąx���uww&�~��Uo՝x�Sy�l�w�Qa��ٳ�����m��I�)�L�=�����M�[f$�{�SX�e;�}��8ɥ�SY����aܲ'kyűFH�88)�Ԯ���W}u����qb��1`�Ccm��R�;�\�1�Vxzr䌨I�� ��X��7�b��[��V �v�����4Jg�J> }��켪��?w�?]�>��{�h���1u��5���]˙�_�������vU<�{J�7���({��P|Թ_|�Sh��I�o-=�gcQU�L�:��h��_#�SP[p�T�~-���xp��NS���7m�i�P���{�g�U�T|j���#���Ym�V^�j�f5z��ӱ2rzO{��\�][� D�s����I	M2f6���N��U�o�Ւ�������:7:��˩�H���gy�!e�n��S�x��چ��Ɩ;h�[�~��xă�B�V�^�z�7V����� �}?��T��ߟ�-B��1���}���W��)�v��q��%��H��]�ލ�����xx[��Y�4����B�MV������GM����[�����f�?�L����g�|=�x��F�m���96�A�s읝�̋���/�V�lr�m
��r�+��]ӆz���pQߟ�?>^����cH�	�+&�e�4V`��v�鰫\ǜ�n�.�veYu�M0ʐ&m������ƻ�Vlu횭*��X0s���뵩��ꛌ�>m��i ڻy�(��sa2���]V!��:Ȕ%B�aF@Q�1��s����w;����c�sb�g��^�*��{��w��)2�%�����Ncl�w? /�x{�ٓ��s���4QI�H���=��� ޢ!}�U�Z �=�+�Ԓ�(8i���7������<<���H�ͳ ��E�RJx�Ɓ����=���$�nI�.�{�8�6�p���d��G�G�*O����nfa<�#ƺT�������`8F	�=b�q��-ԝu�5������a�,�����ٺ��7�p��{�M���A�҂��W�j7�1*mJ]JMD�p�GBN�MۢRɻ����S9�z���w�ؚ`��6�Mc��FJ�%I�&0m�l<�{��g���+��ǂ� ���L��4�rw��b�[�7���d�0�|�/�p[p�V����oΨ���WבS;�, ���d,;��i�P�#���h��{&$�s�S_��=N;��ŷQs���Q�1N��4�D��G{��NA�L,��}3&�q�z� �H�'�$�����uO�߱�y!c[�fU{�J�u���;^���E�j(��#t�S��)��~?vl��]����ka�zi�r']l7Er�Ӈ�w|���$AF��Y�m���F�l3IccL`�`6�~@cz�Ӻ�oX���Ki������U3�6fM�p�Ç�֙G���D7#��F5���� ��ş�m/��O�w�~���3�V\v�5.�u�.�P�K�:t}��&Y`����ᘲ���x xU3�gu|y4�%�J������<�u6~͙���xz@�U���h��fQߡ�M��K��֧>-�T�cD4n���������ܙ1�-����Rn\����W�LP�X�{�\�"�5o;]q3R����p�������>@"P�Q Z(P�cƍ0dجA�1�L�_�֮�~}��>��(�d6`I�*~�����9��6��s2w����L��� ��D���W����6��J{���u|:�,7��>)��?#�������x�J�>��YA�:��/�xx
{�s'y8f,�� %�۰�G�,��~F�W!h��xy��J>�V�e�;��oK������}�y����q����,����G���l�}��V����?�Y��Ϛ����ٕ0"��$��;��Ot�?�ش�{~
��k~%OlG8�Ŧ����F�R^����$h�/�o��M��GCޘqQ�H�	���7\1�6� �^d�F��A��Ԃ�;�q[z.{jߝ��u���OV	�uMִ��l��EY�3��Ցr���J,�W[��&'#3�����|���x@�!w7�k�Ǔ��: Я��ô���l�Ȼ�4/]�y2�a�dVkd�[3.k�����L���^WnA3�k���[�u�8�*�]�hPV���;^��C�t(rl�&��O�%9�q\�	>���`�u*�> �:��X��c���?a5�#�=��x`��_9a��0�ε
���l�ܪ�Im��ܪ�0?Ӵ,��"��D7��[	���zy���ờ(��؈Q���%�{�"PUk"I�qN(��D�
�Z)^��V1�Y{W���zs��;�R�D 8��(i(D7�!0N�TLI(`��ْ9��̩�p�+�0M����6漚��͞n�՝e��d��z�5s��E_V��f�۷sYh�J�ֈ�_��zx7�KC���x��Z�m�Ls�ۏ ��[���x�b�&��[�����l��q$Vk4�9�x5�7i��m�֩�X֚U�0-���Q��TX)%����T���[`�^i���,��j�[0���[Y��l��fѤ�fr��t,����Q.�:z8;��wr��¾^4���,� ��'77�L�0]�@МS��h�ٻ��[��xK�w6/�j����իa��Z�֝t�)\c�������||g�x��j��L##1�ną[B���`ƕ���Ѕ�`�]��6��5��d�����۵6�N�����Gk �SX箯3�*��8u����7������5��R�#('�/e9WU�/������Ls�����j�s$�u���u�<�kͭL�BC-����
,����!u��!�շ]x���vB����ӫkr�ض+�Ƶ#A�رֶ�i�\�i�޺�d�`٪r�����zP���Q�;����M�d�3n
1����#'nQ�F��M�!� ��1:LĖeb����=x�Kw|�'d��r�*���t4�q��Eb�r��^�`���A�W��N3��X�����\ �O@	幋��p��t`O8������wG�=�C��3��,�v7�����=$�|�|�q���eq6w�_^���Y�����H{��b5�s�����-PFP`���Yv��.֒Ê����75�'�+�|�����(H*�r,˔��:HQ�@x@{$�&��4�C���ʀc^�X.&p �R�(��0�h�&�@'$Ss4�b!���V�d��F��	K\
L�[<��ՖD�ܽv�BL�Өq9�	�j��˄��Ҏ(��l�i��=C5��80����E`�n���依_��ӿ?:�=���mX�)��[�;\܄P�UhjhA�^P�s�x�ʽi�s���WS����Q�̵���Ը+mXb�/]����h�F].�9�d�^i�竗��ٻv�2��Vf"l6�ˍ�}wOhb� L�$D&�2&�(43h��,�T��Xy����<�ȶ��P�r���۫�C������|7�qiQXo��'p��y���{�k�+;[��D)�_wU >�{�b�)�L�����l�B�S�z��^3����I��L��7T��:�H��Y���ǽ�2�nJ�G�ah�@�|�-Hϣ�6T������������N�)��}}MVd*鶴�U�Wc�Fl�M�t�s��£��y�������k���� .g��uk�$�,4�rs5�^C��~j��'ro��V��E�H�K�.�M�]t����v������,�M�4$�6���1�����5��z��}�cu�z=����:�Mۥ[�l������xS�v�N�p�A�J)6eo��{�>�'��~5r�G�G����}7t���"�l&�Q��fOx}����j(Ɣ����߯��}�\M���s�cT��PRą������s���C�����������`{�=�	���;�m�����y#I$��r?U7��X��BX�%�p#����{���NY����Yʻ3�M�Z�띇�I���ztP��X��4V���o�2�3�4��6�lm�E��6,Q���mm�$$�%��{�.��i�F[E��7�x{�g�0���S_��G��{����[�1[�J�H�$���?vL�<�#�����DC<���L�F%M�f��]S#3\G蘿5&��a�p�,ߋd�6��s�z�]2#�q2SE��>��x���?�S_��� ����A��B���}_U-8̏|�t�5�L�:��!������<Ͼ�9Ų~ǳ5�1_G�阷?lD��4�sg�&�t@���3�@����AJf\���.5� l{�#�������l察��=���;��)���R?{��{չwd��G:��������b��u�T��n��p�M�4X�t����	򿟛b��d�s��� �F4�~��SM&REU�/�� �t�ʟ��qv����� .\��$�,��[�bLaK|��u�]�<�#T�6�MۥZ=�����'�gn�gG��4 'z�f�2�E&̣_d̞ w��I�?�S��ɕ�q?��UFY���i��nQ�T�YK;?c�g�~
}g}2���\���9��V��i��(J��-��R�p�4s�*F9�(h�v�՘�L���nm�n��)u�]���	kT�[��su���K��,<n:�ճ��c�7S��Vg\��9�}s�V�6�&(زA��c὎����g@\Ⰾ�y�d뗻�����2ƍW�����?��bLU����w�3'>�e��I����<�c]�fU{�J�g �B�f��������1�"�w�@��-E�;ӎ���%��<</����L�6�_9��
  Xe�vP�.��F���$�7�^�ʒ���WPzJ6m�(�OP��5̐�QR�إ���I�ɂG	-ɪ�n9O5wS��:� ���gW"���o&�	�J�ټ��3g�X�C���#E9[Nj�h��ϑQ���v�>�:m�2Y���6?���c�01�1�E& ����5%o^�1Z�Σ�I+Ξ*��4�eG>�'�������͵?il�Q}��S��B��xxy���rw�d������fU>��l(%�K�^'3����j��%{Z�1\������᪺����<<�e����i��nC���S��li��p )|s�HϢ>R�%K?k{�xS�ۙ47��&0� ����be4���'�i��l�`��R+g�=�&�t��WDV���*	��������h���.\Y#�Ȕ�a��z�M���2���e�
I��G�ޚ�cM������ od�j���2�%�j���W %�w]��rfM�p��)�8�x�휪i�a�v��q��v�E��e��J&ͣ��̓��?��z������gu�"\'	�T~ݟ����1&4�~���`��ވe��I�����m����U3��̚��қA�3.����Q�ٛ����`n�NAP^�LO�=���̨����'�87���=���\���/�Pe�Y�����)1y��������{ۻwo�ϼ�{�}��\��5j�k]Y�)��m\K���ھ�ڰC�ܮ.�}�����턣��pnm��^�������V�Fq�<̏�����4����X=p>��n7C�7m�5�I�:=�}�]�w��w*w�G�j��{��E8F!]���~���55$~����P0�D��=v���R����h*;S��]$C��F-�
!K�g]d���1�����c���Nw)Ƶa�׉��6�j�H���֕K�qk����k[���y�H
h�Y�8.�Mn:�c>�H�[2n�l��	����v�ͽr���u�Y(f��:��^��s[��8��Y�㇏��w�w;�:w�C������ɢ�x~/��'���T�ch���{ p����d���ICH�PԾ�����I�a7s�}Q��m��*G��Y�S�����cR�����L�YEUX��I�t�ʟ��Z<5�U3k�&Y`����g���̣��̓��;�-}adCQ���,6�V��4�+��./�A����-�Y�sh����O� g��O����i��i�?f��6�SY�C����x��n{NP-^���0m&�ġ82������Ɔy��t�]�/�I�\D�ߵU�;���{��1Z���"�̣��̚ވe��Ow���Okl�������۹5�>�i����G��o.�F���Bw޿��%�	�JmR1�f: $�mZB
;[w�	�L4�ܟ�m�����Ͻ�Q��m�vZmTO#�ÀSs�\��[g����
J���Xrw�����wR'�CO�{��Y�s����sϴ:�.�cJ�Kq�jj�\��C���v���!�5$x�����c6�!Dxxǉb��0ev���(�j:�fk�c��\��d��*;������-Q�dR���g
���-�=�[O�=ow!9��%��z����%�Fz�^���=��/�\������0m��cʉ�{��Ӈ�Ç}Ȅw
<��j��/7�N<�9�r�{���w�iOa��/,��)9�;ޫ&�|'�eњ�|�{��+�-��~O@�}V{�eߑ�E��2��X�;�e���Q#�^�4�]:��le��w7�i�is]h!��[��#]D��Յ0#��w=r��Mc��[
�s�:�NG>�b=�s�c�Tp�9.��]ukͅ���8d����n0E<�4%t��,l�԰�E��oH�Kl����+�'� ��Ź#�j��#������`ݲ +B�c�&.��j�`2ʇ�;P�M�N��
q
"��x����� Q3��uk;O�nz3�d��{^E�L��̘2#�m�:mJ���{��)x��Y>�;�<4�hlꭒ��u�Y�%�ǚ�i���*���9"��
�k���(���B��p�����=�ހc���J\�CԳ ��5y��f�`��D/!R])��$&E',̊����}��sVv��A �f)��T�+<W�����9�8�	/C��9w��}5��%4����,aӢ�A���{8<,��z��23����ԍ�n�l�[�G� ��{[��Wn5�x����N��H��Q�Iύ�Q��Q��FA���Ƿ�N#阻M�l&�Hu��4w]Q�m���t�{i��D��C0�}��'G�x>�~;���-���3��(~!��(h&]b�y��؊��{W����9�10���"M�pů����mT���8��$�����Mnd���]���mr��i��Kj����\���Dxe���<weMG�#)��H�+��<�2�^m��A/���ۀ+}�����������5�uY�Ƞ���x�v))x�^���pv�@Ʉ��y��|�}�e�UQ<�#��,�Up�9m��ݿ��}�nN�z��-.��^Hݢ;<�W(~Q���
����b�G��8]���7��I��-�Up���ov�=���,�< �Y����e8NY��d�1�|o�SV[&�$�-�U�_o|n����m���uRov!�P21'�*{�['��w�fK�B��)�WpV���L�UK'��wr����,_E<W�a��2Hx�v;����%\�O��]g���tC�͠�F�,s��\s�u؉8��^����ѵ�N�,��+7���1Ѩ�h�ѹ�����TUqb�v�n��ı��+t���֐���h��:[-�/2#�ܼw:��]�uӌp��[2�Y���]�������CzN�[9W3$�? >R�;����7��2O����2�Nj�I�xހ%v���p�h�Tm|�2�fR���^��%����-Ώ-ޚ����\��	s0�|�f&���Wal��۵R{2fM�p��e�1����i�j �����)�. �ֺ3T	%�=�3$�0���s}��o����n� ���cs�\�z��p�1���#LE
�5y����P�5�%�Z��50^�t����wѧs=���mLm�#�>u�]9����,���������I�?���[=�ٖ{2f~\���2�$��g����S=�3$������wB*S(�������y���[�~|�)������|��N�c%���4Cd�K�4q_׽=�t2��'��l�ʞ��ޔ�[f���P�	$�ާ��TaH�\�Ԗ��zT�����a�*�-�9�*rψ���SgF���XhC����-w��ؓ�5�o�z������~�y��%4	��� ��ׂd�'�ْ�L�ɕ��''Q�~7r�|���s:I��]Q϶z�| �scJE�l��;��4!�v��&�m���j.&�M$�C(�Xl��\�$O[����fM�|�a�n��i\SR�:�#�8%WDp��A�F��m����z�j�f0�v��(a�`�g�����K�����OĹx����LH��(�Ѷ��{�6vvB3�cGf��ֳ�ieLۈЙ�I�<�Ͻu����7�&�8|<�r�[l�@�6��~x����7U�ձq�t�8��.�P�+P�]m�}~~4�u��Y�èD�7�Ch���W����0�}�3P��k���S�I�1
���LɽN>��]ZQ8��A��I�����seGZR�uˌ9�Re��m
�7��ޫn0�����ۑ1�\IJ�B(B�k�Gb��Ō�Zl_IF�Ӎ��_�~��2�V��r��n3�n�Ǝ��f��s�m��,ۮ�F�sn���c�Srv��J�F�z���;y)�	c�-��Ҩ&Y�a ��m8��ٖ:ĜU���]!�M����!��[e��,�z�l���k��r�es�e��z���\Ŏ����gNqM2�Tg%&����5�<"v3Z��ڤ��j�}���cbw2�� �y��mAa$���ᘫM缪�Y8�����&S��=�E�J7�����+�g�e4�l�5iF�\}�l����{���6Vw=��#<K�(�� �ڂÂu}��Z��xK�J2�0�@�l�okڭ�˙#�_I�UQ8�ˉ�ST�@��u&C��꒑U�����{fs����u\�Lbm6����lm6؛;��[�n�7����z]<�L4>37c�W2��g�=J���?n�������Ԟ��f�&dާE�K���M0�$���< s3�['5�S���'���/B��5��)[�F�S���:h�������|	���3OG��:�#ƣ�m��dҭ�ޏ%�-�왓z���;9��(�h�)���R�br�Ξl*����IA��J�S�pv35��q��j���Uv���|�|���]�������G��z��l�U��I�L*������Nr�L��M���w�L��K�!8D���6�xV)�w�ٞ��9�{��Ћ�d�v��tX
�\�P܆Қ�M���m���?�??U/��ů��Xt���I'�}3���{�2s��b�<`
��Ev2�a��F�o<'��TN�lҧ�-�XI': Y�a��M����tET��\���l�uw)���	̭�0DH����N�K�/�l�޼��x��~�t����h7�D@��#5��L�f�\ch��͙�]�2~�s����D'�"�@!q�՜ݺ��y�ة6qD7wJKb7�B�4�'�����y��E��K��$�jl�W3����G�[f$�6�-���L�]�2ky�u4�_���x#�)g�&d������e��F�����xxVeU�ᘫM��ܡ�r�.�X��^�F���n9\�z�	�Z��g�������Pu����׋)����sl�B+�g]�2)Qa�*5��1���Y>�}�ͷ��3� �F|�5=�Q;���F��%ֵ�F�fU<�k'p�⡐aΦά��XJ`m�c1�=�w��bk~ �U���9G�!�U��R�;�M�E>��PĪu&�/��t�Q]��&�ˮ,�������"f�>W��_m����v�q����q{5A�k�����l���=�����I��'��잡L���C����Bl��)�3F*LD�bg�w���.��=pgf�աwCcT�C� ��kb7���(j7��3;�s�1��[��I���r�]�P��Ѝ����C��5��[��.����r;'�zw���M���彑s:7krNT���ݝ�h%TF���p��p^�u�+0]��� Àx�ﯯ�>�~�0��� ���]��oc�s͎{������-�N�=������Wc����4<��͹��8��k����cM��b�iYAɃvS3��|e-$���t�۞ӹO4<q��u��O\`VS˘Ī�U���ڃ=�z�X��[g����:�]���$Ga��<ٌ��6�xzD���Y�ݵ����n����w^�랞�Kj�u�1g�l!����^q�\>,Cd�ۋ�����L�&��N�F�ԛ��X�T���\dو;P1f2�t�<,ٮHcs؅��$e��ە������	���u�Ժ��'��cPu�KgY��Z9w6��Y͐�u�6�t݁��n���D4gpAۥ^��3i�`*�B7[.ȗ3Pm��*��c\�IV#]���l�;�T�̺�A6��Rז�.�����3B[jcKu*`�e%jAWZrj�P��^G��.:���2�\��q-ā�V�#��Ԩ���i`��՘��-�x�YY]��x���XeQ��z{OQ����պ5��ù�úm띢s⛝Ɔ���rڮ-�b��:���C��&2�N�:5�D��Tؠ����&�#T��#pŪ�[^,��~��R�;���C��n�	S|�#;���@왪�3�M��������\w��c��N��2͔j>{�p/n�(���0���T��~6�~�;�77�����Jf����W�$��>�a�8������|A��a1����Zi����iG�5�̳��s���D����N�ڰ��ժ�,���^�3���{&��B���wI���`�v���挓�o��p��lIS�/c��Y��]�z-!��=Jp�j;�vnh��F f��U�"��=�HB�$!��h�ڝ��-# c���y,&z����l�ݭ-I��=�������m�8�]�b�ٹ��cH]����d$u�÷��k�m����F/Q��&���<����wx��
�)�l@�+��YwNF���=H��Uf�չ%��%ޞZ�3��UW�R����m�p�T��+��0�X��`��f��ד2O#� �?#��[m*u����ޏ	U�_U-���*7��Q��J��y}�U$�0��s3����F��Z�BP�UW��p;&d��,��̜�o�Ϗ�[W/\�[!��sKnk:m]����:�s�7*|����Q�����*�&d��C�e��?Y���G}�k��9�ؙ���"�K{Zf���Ŏ�"�ᨆ�����ӛ�5�U\��sH���SAM6�m{g.]���3��<<*���U�#u�f�g</��D��Y2����(��0j��/��s2fj5��-ٖm[�[��NO��b{��2�[l�F�*��\�n {>ۊ�ԼGc��%��i2�"���kh�6���
���<ÆK��m9f���#�d���x J�j5C�!'Tw�fM��M*��ev��dG%eg��`�4�:Bv�9��d��Y�L�\Y�� ��F��F�ŏ7�z��?<�x�9q�@�l��������{����U&��94�_��cy�~�yUD����&g��!ѥ��HC,��IE�Ab�VPݥ�V�Er1���?sl��̟�� (��m��v0�������̙���N�{�J_+��p�p��Ѽ�$^6�{ʮe���<f>���J�k �,���޹���S�Tn�M&rv�b{�7�Է^D;8>s�\G���q��߮��h؈Ř��B7>u����=sﾻ�(�0\�x�:<��g�ə�J� 	3���$�gk����U���l�ɶ�N!(f+����RY�bL^/�+�ə<��A��I�?n�x
��l�����=T��.I����qf;��ڹ�����1�g�5��Ҋ��=�}U'7fd�'����~;jl4��'��r��w��;m���\QMߨ��)ƵL�h�/!�a= ���Hӗ3��[�;�����(j!���L8L��P&ձͤkn�u��sH۝�x��.��.Մ���Y�k�����j�l=o/�=���y���.,lX���F���[Q3��nah�;2˰S&X�)Tf(Q���w]k��(#A��hcc`�x��uvF]Y%��1��¦㛪�VIv�u�I.�_<sb�6z�xp�I�a�g��ni�up���fKg�ə7����GC��-�,��3$�0���Sn㝄��tay�Su���7�9�*/�Us,��q��I��e�x-���=��d�po[,�
a��%0�A*\k7�{8-��{�D}��4۴�g�xR��˓����PN�w[9�������wi���&ã�q����P��0�4�7��~��>9�����B�1Fd��@6'�Q�I\��)�W8fgg8��P�UD�8CQy���(�J#���p�0\��/��L�nJ�J��]�Q?+X�"�iB���@�d��J'!}=����dk�b�t�)�!��p�L��a�Yi*[���e���ri�V؄��0�:�xy���c]V���gu�)��n�������T^f�s�s"e�n�/�����_|���׿�9�6�,i,llʱ��Q����{맞|�PT4�� q��b����ʩ��%!(���{�s2oS�cm(�=��g��:���Vrl�W���u���E�m��7}"��k�=2�[f�t��L"\����������̞+}��U��m�YF��[g1������k����P�M"�K@?f��1��̪���3M���g��LgGw���x�!�ot�d�ԳӼ�\�i�I1����)��4oWWLb��A�U�ݙg���QF>�H�[w{�a�O�ѡfh8�,A%�b�ef��@nf�Ͷ��"��wL�cl�> H�V�Vh�Za�n�#�>���2x�G��=�����pș=ͳ4�	W�a��j�O���-�!�N���8G3.��r<�Q��
p�0Z�z�=��7�������B4z�_ӂ1�}��\�$��*=�ʏC�������2&u�x׍m,�i٫���i����j-��W� p�¾6�[�rV�);v�ͦ�M�\����Ƥ������5��9խ�k�cŵ�Ĭ)+r⭎�xb�ūkuƮk��������ۭq�s�{��pL�#b�I�%F$ڋh�
*,��b�����;��7{��t:���N�a{v����v��f��Ԣ�(���7�F�g�0�h���r�g}��=�H��#[�7V�{�k�Z؄�0��kl�'<%Gإ������a�ل�DN���uT�H�����e��5q�PT4�ѵrl��ͪ�~����1��}����nv���m�nQe��نhTDWD>��g?y*������jl��~l$UD���f���G���/zG���sÞ;�tA�4oJs���c����c�" �cTRj4X�j(�#&�$M@	b7�"�Y�WUU�#vޏzUw3M0�$���X��Ώy��U&�3�[�&�e�QSZ6�c���ۑ��˿��	��-�9+�jd�k0�fL�V�9������u�Zd���X�^i�%��h5��N����^Lɏ�|<$N?�j�������bO۳���G��z��L��Ɩ�jI��Yʹ�5�c����ד���[����UI�i�ו\�^��P��1ǅ�������r2{��n�p�|P!��c��<��xLV������8����%�xu@���=�.Oh⇺=�3�_��g�OIkyW����ݏ��{���o��Lzxe���P�#b0"�䑲 ���frZ�!׫2���\B�q��ڗsIޠ��;��.sW��ى�f��*�SKk��K��mHʣ,ƪ��~���vq�~�er�?�R/;�6�4��b�6�%��mi:`⑨�ɛy�+3}靈v�9����l��9Տ�[�;��w���mX�!��*Rgwm�F2��,��~pw��o�[�~��=��hwZ��"n��zV����{ݓ}S�r8IW��|��M�h˝˚d�Oqp�=�h��Y�nNY�G�t�Vֲ���N<�ד�/^Ӭ�TNiE[��!��ʵɹ;� ��ɲi�"N�:�=m�[�o8m�T}t'�fV��վ���X�����~Y�f#��[��y�FG�+O?8�|���n]�rd��R�~i���my΄����}�'R��4��agoj΍��F>���O)�*��s���>n�3����ޜ�7�Tt��z��z�C�z��b�t���y�M��ٝ���i����+!�R*�܂��d�p,?{؄I�v�����`�*�r>��j���O���Q�ꯌ����b4�/E[��@��b`^� ���v�۽ⶅ��b�ӻ�� �%�~�ǯ]m�mF#!4Rm&�TfF�J����X��nfOi('/����Z�缯Z����p��p�'T~=�=��?bQ֔g��-?�$!A��s�q$0WZ���sۖ�N�	�Uݾ�Z<0��C�7	&SJ]�����JmX�T{pSf$��͙�q�<�fT͓�m[b�` �Xv��_1�9=wY��:{TV:󈬚%ïj�7+5�`병�c���q�?~�}QI6"�2IQ��(�"!��i�cq�N�;��
�N�;�_E'���^�VB�y��	h��D2���`�iSO���A2�����7�C^ϐ��=�Z�0��=]���uX2��z�<��kY�FF��r����u��0�f�ݞ��!wuxZh�-���E25l��n,���[h�h�3%��j{حK��n��2�0�ia�km\��a���o1e�,�D�;��S#V�jm��K�R\�-3i�r��h��=�0�k��b2̵l�ia�k�{>U���#���x���y��E<89���-3���o�^dn�=�sGJ��-�]M��d1KgK��J���o[,���1��jz؎9ۺ�jK�Qsj�kf;X���H1��[�RZ���z�ض����[roq�^��hu�$�ƝΚ�fz�\�����ǻ�I�hѲEF"�� q��8��v���2I�OS�t3+v��0vM[s4R۹�˩uRK��l���Z2�j�*�L�[+��<,֙���r��h�h�9�u%]��-4i�׽ܸ��ti�k,�;k,�Yh��.k�k��,�CZdk���IXE3-[+��Yf�F������,4F[\���e�f���ΥB[�ZfZג�K��k�-e�~���Πj��E�a�G�;Ue��e�Mr�e>��ޭk/l��0�5����ᆰ�l൏z��6��ݪ����n��K���x�j��ƾ}�{��Ƿ��rt{��qe�k-�pR�Df�l�����p�5
|
�� 8�Yà��"�j��m:��nRS�3ņ]����5�+jD�,<�]:W%��r��&hj12J@Li��hl~���nk�뙋-g%)�U��Ff�\�H컕d���0֚9�Y���lܥu!ᑯkz��2ճޥ�a�4;�ow#�rT�������Q�{��Zh�-��E25l�kqe�k,��l�Yh�vs���n)���dk��2̵o�1^�-3Mi�뜸a�4[=��,�e��R�|�ˠnu����vC��ʺ���#ku��X������c�����'|����a�2�Ը�Xh�0�w��e�j�+�}��]K�-25�������Dgw�E���ڿJ�S#V���Y����׫�w�����E�ڶ�e���?
�7*�K�N+J�$}����C+��b	4�G���n�QZ�/�;Y�)�F3E##14i�/�M�|ﾷ�ư�u�\0�-��9��H]�Y���tE��U���W7Ȳ�5��J#Q���#Q��mc��f\��ww�a�j���a�kq/1j�㽸m�4[=��,��'c��w�:�}�����������:�URB�f��\����t�Uʔ�+l�[h�5-�մ[-�{9��8{�u�kL�ia�k�⫲�R]���-��,:�4g�hm/kv�H�nѴ�)��{�u%]�a��s����i[�e{{�!�����KZ�ͻvY�0��>������,vY���u�wmQ2iRܳ�S�>���}��8h�V,�޽�O�nT�h,Ңf"��3FLcm���^\�Z�5����T"�3G��Ȩ�? >ީ�ł 8�׊`L	?];����W��4",mA��)l���8��u��ۮ�v���2����0�0�x��a�\�.`S+��d�r���S\��^C-�h�;~� ��c��(軄��'�%E_�=W.7PC�m�E8L���={."#�n|=X��)�M�RSx�o�������R�K�v{�)RюVG�.�,}%dxl0���mO���'?no�����������1���&����4M�����ڛ��F��l]�n!��]��14���l���f���#WF�Mp-�[��+e[��c���6���Q^�F��] K��B� �΅�#����5���e�T2f �F���w�b���O8����kvW���j�`�}�?_���Ǻ:;������Y�-��1 �)�����n�p��	�-�ma�	偮����n�e5;�F��FX��>W��K���F{��a�L����P��k�Hl���v��0|~)Pj�Q���j�]U}���0|�5\��ߍ�	"�����-�A:ޭa����#���-�֑�|���s����]4[5���"h�ֳ]���=g�㽥���3��!��i��G� (�_l�[F�ܖ>��麌 �v&Ԝ��mLKc�\�#��qK<o{�����S���|����Cbn4RF4V,_�|^�]{�a;@wt�#�K{�j�.Yu%�6{���UHo���Z��݈l�5ݻ�*�� � �-oݴe�b�)FF{[�a���*3��e5�sun��ٖ��Z��^��a�L���js6�3Z���$.S�G$ue���nŝb6����WE����A�{��!��݁��ttMS#GuJ24t��V\r�e�h�nW�-�kV�4��V�>�W��4[-{�쐩R;�,��t��h�iFFo�8���ڠK��}�8��왇JG2&�N�HŎ&�l�������5�!a���͋Z��lBm �+�q�L���j��΋��"�f_R{���0+���
g��@03�.�%!����܍܅K�,�vY���@FSX��f;�Q���5���]EA#R�� d�w`��S�[M�M�RT. �w� 
�cک�ѝj�!�i{���o��|����2a�^��!�a���	T��p���o�Ymw���AՎ��̴{޵�a��K#�-���SS���y���];�e�����޶<"=x}�s�r�`�l�P�u)�}�c��/S�6F����u7�{Aan���w�ב�ElY-lE��=wּ��{^�캑�e0)�o��.RV��]�o|��5׾y�YD��r�����]�n�	B]ˋ�X��Tp���;@���Kݣ�ꂽo�y��U�.��Hh9�r����h�P��˴����%\�WXYzh7�bA:h�H���Q�Ͻ*�.Yu%� �L�w��#F���mF���y-'��}����R�F�H�.-�w�b�b}�Ǆ@�� q�V(�����36�����⨩{ˀ��k0�Fqo��cQ�+s��7�Q9��,Յ�(b0*�s��L��$3�b��<��:�#���u�A�q��R.g�^5�m�w�&ʎvr�.b6[Jl¼㡕*�Ex7?K��0%��Sz�p.R�{�����ox��Ѻ
;��2�͵@�b���������q�P65��/*/��0؂	����N���Z�B�`<G�k���y�����7�3�l�!`��\�m�aν�8�\�M�2�^Ef���4��J$�=9z�8�ˇ?=�ƈ�+b�U6$��o��>��*��Ԋa1B���d�0@ۘ�[���4�`��S�(u��b��k�;-Z���U��Z'6h;��*E��=���e���r� ��7o9s�vE��� >s��gl����=���Ɉ���Y��1����8���!e�#׃Dt�5�-��$���5Q�L�IY���'Ppݺ��uʺ�T�5٪t˶���M�i�n����5�v���G%�:kA�*X��s��:�N�P6��7>l��H�J���� �u�Ktv��CW5ĳUc.�4��f��\���jXF�z�ݚ�:������ĀE�Z&��F�[��Eź�I 9 2�%��Y�Z�Y��@�-� �+��h�S�"�c�)u�9�ƹ��Qr<���t]hK��EC-̺�c\�\V��#��ъi��x=Q�\�J��\���Es]^f�r]4Ś�έL*�M�udՎ(qۢ�fj�x�I���k�iWK�Gg6�SuأWRl�t�ɔjl;B]�s�R�pmڽ^�[�r�]`T\�y�+,m$(dƹX.#4�͈��� lsκ��=� ��]��y[�.�K���k�bY[��6=��vk��Mٺ��"b��ɮ2�.u����ۜ
LlV/�,6Ҵ�0]����/v=���
!b[i��g.���:��7V���F8�G>ql )۱�o=�涶��r�u�1�Z`�Z��&I�7�ɘpV����5�+�0G��/x���2���#�rv�iwoǍy�C%����32l�Q�{_[�8��䛷4;5���>�g��|���V�;C07������e�j�vr>��$F���,Q��r��U{���>S�� ��tH4�<^;�}��$SѦ}���ճ�<���C��� �;$� �#Yf�6iH)�4�^#d<I�.#C�M�	iŨ:��J����,�tl3UNT������2���W5��$��y�v��sb�v&�l|x�X��`c��%����/��]�:�W7��^DV���5яC9!!KJ	i':T�a�X5-�k�\8:Q�s6���ڐ�9���oZ��)b4�ۡX1q1Ri`TH����ڂ��t�+�-�i����hИ����@��c�<�v�y%���t�4ڑ��B����zN�tM���ěBA%b�QU廲U�&�ҷ>�F�fl���Ү��n�����j1�؆̳�1[D�"�X·�¯-e�A]�n/iS;�X�uHm.�6�4�p��.9X��4\�[И��Z���\ُ{��*Gx=AH雷���ڌX�����6�h����΋�"4S;�Z�F�]�)��-a�N�M͂�s���]EL�X�F���[��[BS�E���HT���F�=�h��5m�1,�Ma����F�ђ��۹\�*����
f�T`��r�)��./n*k�8�#9[F�D��tE�at�Nf�֮;�h�k�Ԯ>� e�lmllݍklm��5�k�q~z����7�h�R-���}������F�9�h�ѭҌ:���۸�»��h��^�X�m��e���a�|���L�V�lؚ�qh�E5���v�����Zb�EW�q���i�ov�і���E�[;�Z�F6���ҥ���m���jn ef�;C����ի��^�����ޛ��J���h���"4S;��}�S����F�*�.���l޵kh�e�4S9�Q�@�5��u{n�UXF)���<	�O��f������J: �;O~���=��{?r��8f;bM�릆����6r�c�2�Ia��I�@�I�&��&����]h�ES�j��g�8�L������x�wJ��07O�4�Г���Xh�צ*�]Gn������n�0�v�)���f�0��KDh�mѿs��:!cn[�UNXˇfz���cF�:�;�im�m�F�f�J4F��U�K������0Ѿ�Uջ�t��h�s����2ѽ��)��(�1�h�1H�d���W�4�U�[E3Yͬ0�Y���E4S7�Z�F+g�y�Q��0�[;�Xh�ԴT�[9�Z�xL�������^�,��e3���.�ȭQyO�d�=�v]���v���^��=��yכֿ�U+X�����amS3�{��R�w��i��uh��~�|�-a�M��F�guJ4F���{��gĨ��Xlh��]X��+m�b�[I���]�7Ϻ=�o���F*������vt�FZ+�V�a���9$uR.�Ѧ�vZ虆�gZ��h�e�4S1���6.�Zhsu��%\��wxDi{����Ջ�0�w{���4k��is���F�ۅae��=��l�hh�kQ�b��kGk\�H;���V6{��#]���b�T�w�Cfy���ˬ>b��nL��s��8w�4�x�9��Zr$����ˡV�v���)O��.��$h�
P�&�c�˗iR�����֤�%�׵�nA�Зm�s ��V'�tI����ώ]u��]bn�+��e.�[���h���cՠ����/�=V�]�ЋM �e���Kz�v�]��\�O5�Ѩ�"5�=���w���|���I�i�+�e�!t�.����ֵ��0��V]J�h�w���yq�~�Y�A�J��r���}�UJ�"�^j���k�ٶ4n���#ť�u��$�uu��!��h��f��Xa�-�-���R��>.]h�
��#my��ε��h���-����`lMV�o�rUʕu�e�ݤ[]��Q��u"�;�[Fг��y���R�
n��N������מ�i�v�Z��I�[���=:��Ρ�w���%��j@q�>�^���߲����LH�;n�n&^�ښ#7�i�ݥB���L�滌�����/
��6��lm m$؏$K�,�y���Z89�*���u�]�mF#Ԃ�0�[;��3��#K�{�*Ʌ���4W��Ll��`F��!����wZ������Y,���t[����H]�u��{���}��v�=�3=:�<dJͅ��4:ծf������ܳ�ڌG�vtC�nҶ�z���!p���s�@�o�����X��H�#�_f4���iO�n�>��QJi������`����45GN^,�o��]P�.���a�_a�|�CT�]\����� 3ș�C�զMR�{�j�f�ḳ��n!(�O_h��5�^�X=F�q�����6SUͺ�I��6@�@m���C(��ǛO�-���3u�-#�ѽ��[x��F�_��'#�$���U*�=^�Fi���8�)�����Q�ݤ[V}y���s��x�p�Uk�t�î\�\Thu�mv39;��Z���g�J����h^Z�-�������5����g/|�����Q�zt!�b1̿U��rE�9�on�AWe#���1ld�[e2�4 ������z�������ģF��7r�RL"�^�-G�+n�l��`F��JK9��u.\$�,��dٝ����r"�^�-F#9����x�2���Ҍ9�E��[Khk�� �����p�$�h�w�-� }�-a���Cgs�4`��pU�C(L�_Nj{��"�F��;��sS#�E��z.��,,&.p4a�ua��F�L&�~�������l���mb.�A������ۧ�c���[z�`OFb��2g���S�"�Y�%�v�R�a��S��f�c�2�i�����x��ҵ�MkVwݖ�IoN��=�����e�n�ʔ�]%�I%�:�n�,�O�0��z��:��X��E0�>q&,4f�ȋid�ý�
%H��b.�J��j��^�"�\�+f�0+��ˎ-��e5�z����V�6�/o���=�An�\~֥�Wr�]��T�v�\�+b=�ȃB3[���K�U˩WxE���Z���ۤ��_y�`mY�o��l�˹UQ��=n�z�9���{hjv�n�n��i��; ���H-�խC��Is~��#��_$��B7���,� &sgЎ��{��^3���aᶗ؂��ɨ�Ko��r���,M�ь���;�w\�I�<ы�[Kz�lF���4SG7�v�˩���2����-��r�aԘ�n�6wZ�#C��UU.��k�a�ҌF�6s���Mr�~
=ﳴ��e R�Tء<32lSG�Dj.�ZO�{ƨ��dmպ��� sJ���f�����%ʻ�v�Wi�[[����܇A4�|�hѫ�nJ�R���0=�-�A����uiF���H�:���˒�I0e��; �ֶ�[�7^�)���|�j<���ʰT:H�ͱ���V���׳<���Vh�8���I�m[��q `�����<v_ ��R6�ͻ����]���Cd��BV5�&��v�`�`�q�_�'�����x���8"�D�W\��}��-���W��9�	刹�F�t�V�Ҟb#N�e�j��5�X�v��s#
螽W띕qoV��*�cp��u'<�*9�Ky{�}���-����&1&�;fR�����~&���=�L��;A����-ў�A�/E"����^��a����PU�bF֌�%�!���l�q��10��ĕ�u`�D����)û2Ţ'4�ٚ�Enc�,�OD���wGR	(^��V7���4g�3m�MH��蹗Fzy�q�wz�f��ˌӯz�j����.R��q�Ӫ�d��=�C6�1�z%vfD���?�R{����)r6oҟ�Gbg���=��/�s_m�-a��Zц�$;�x�TO�=���e��W5-"��ֽ^�1K���2�UlB.��#7D�n��({!p����Öl�ϋ�'-���z�7Nǔ�3B�sP����	�*'}����Ou�C��,RZR��]'�˂��	�@J�8ظgp4&��?{[�C��ɯa�c�^�o����;� ^[�\K57�ىӿv�=�2�΁?lBa�B�:]X<�.��ѧ�lU}BQ'9͐��uf� ������f����+QP'6�8�
�J�,`/۹����pl�������0M��]�Yf��F�F�Dj4����K�	.adq��֨�^��
f�-����ᆣ k��b�J���u�����%����mky�(�Xi{���u#6#Z��յp%�n��i�e�4��Žiy7ѹ�_>������05�oa�Mn��j���;7h�Xh�Ύy�K!�-e���Q���n��a�5}���h�op�\A�:J�����J����J���V�=kW�m��F�.�Z�*j��Z�q�庘x$�shmF�n��j4��b6a�����x���q��^�wC�j����%y޼���������W�3�ҍS+^�$��ܻ��-��o�F�RO|Ŭ4��kx�a�f�-���={����J���(W��$6�n4]h���Z���=�z=���ߋ�������0.��=���8�q��R��� ì����w1`j���|�6F��c+�r��!�\�R"���Ǧ<+Hq00�&.�6��������T·��՗R���EH����Q���a�M{�Ҍ�ٽ�0�h|�j�UR�Z�.�Z�*~BǬ��ؖڶ�t�յ�Ʊm��3o:�8�1���K�W���hN50m	��նpg''k �'�[I!�L&�Kkq���&X��jm5Vv�.��F��=z��w��V����8.�M�ۦ]�G����v>5��t:���\�eݻ--۞s���M�zH7oGg\��c�\tGO=1n���s�%��DFɢ��ÿ^3��������l�R�[�t�iL�W�������ݯ|�}G��z�:>�Xiwr�iSY����.]V�T�t�h�op�Q��sa�Mw����V�nz�%\�xF�G;Dj4��j0�յ�bҍSZ�Cj�1]�%�$�2�kba�w1e�Mw�ҍS4�m[6���5��y�v�]�I&_���!�%Z��\�"6���Ӯ�s��=[����G�[�c:-�����D6s��c4�is�u{yb5����Wk�tU��2���O���q����6~Uk�+"r�oXKX�[�ne��+!\�϶'a���g����ߍ��Ũ�7�,Cf��G@k�N2�d�0��[1v-�aLϨh|բ�[ǵ�J�w��� kL�ZQ�f�H�F����a�s����5]�r�R8\�S	e�e46��foZ�Z�I{��YiS�!Pg{��'1Ƒpu�RAkL��	�[V��e��O�������3|{2�e46����z�W-ʫx2�i{~�>��mw�-(�3{�F�FyDkib��1^�Iuwu
s-*k|����"=8��W1ק����2����1P��Q��z�y��Kl�'�}{��#�lM��=m�Hm$�,4���,4��^�}�uc�;0�_�2���0�h�)��[K���e�l5�o�]��o oT�פE�x{�Xiq�v�j��R#Q�`WtΜl��wd�w���qK�����m�Fw�}5]��T��D��3WGj���ox�{ҫ��Iwwx~�R�ot��h�h�F�;-FqE����WW���3�Bm[F�Z��`^�3ZT�{iF����nJ�R���ĊG;F�K|��=���_�0%nEfQ��7wj9�+���.�
��t#KA==u\�f�tBɎY�s�� ��RV�+�*��n��2�K��"�+������������������N���ŋa��ӓi�*u�uu|�������%���]!�m��K4��﹈�Ҧ���n��.]�K-S9��xk���泌Ҧ��b#i3-[5ޮ��tU��k-��j4���,0膭�w��ot��h�:ۛq®�����0�k*k;�"Xj���V͠k���,#J��U��J����J��ab��orc]��K���t�+u0j:���sʘFrk/Z�r���젴K�Ja��oC�<͍]�;��;��\&#l5��ַo\�Pw��p�+;E�HK۝�=u���ַ�Du�I���=��\f�筙 �ulܛ=�.?jn�=j8�Rl����XG�w9k5����c��C�gf��2@�3\��~^���u���yoļ��1Tn��\W���s,f��8����x��:[��Ρ��K��!��Ҷ��ZQ�eg��K�Wr]Vme�}�>�f[�-Fj�Ϸ���n�H�Qᇮ����\��Ȩ�{�\��s��@�S{�D�7���I�L9�����01�����od�F��[�(C�bZ �o~JSq�������?���v�l�POn��nl�\%j��-Lߋ�>�����k��{�3v�݋��+~K�Α#��Q]5���Ղ'Y�$����#�{&8^NL���L�	ݼ���������s���v��w�N�I%1� ��g���AOP�6�)��9e��k���<wXQV��e2�9�Ho� �n'���Ag�~�c�,Ge=4;]m�+�͍i�V�-���u�������o�>?=�u�Ee���ICnb���o]�u[x�^��(�����Ue�_\���v��=5"��n�6�A��������W]�Um0�=��e��[ 5���Dz��^���e�w��ϼ۾8�VLUv�=�ܙ��|s%O����`�AP�۳S�G[������n9i6S0�a*��(����oq(�X��e�4�6<�c5�ģmg�Q�Q[��E&�ID׽�<>ߞ�_�����^���/57����w�3�>���x0���6�(Vq�n7aM�Φ�콪���\�Nj3�(#6�R�U����}���)��}�5u������S�~��}���^5T�X ��� ?0Y��H�f�]s�R5��\W,��!���n�[�~uZ����%�
'�5����q�R=w#�#w�h-%/�(���t�-�ƺ�����)Ow��P1wmΥ~�cqZ9�8mTƜ����]��N�bu�&����~�S�BiP�ߋ��O�:҉��滃�Ǹ�cau�UH~���T���S�n�m���ᫍ':I�}�vW�/xv��u�N�GZe�n�٥ڍD��۫�B�[/%%%^��E^���H2+^�3
�����U�	u���Y�{CU:��E-�7�lq�$Z1}
�Ѩʾ��T��˨�x`23��@��x����~�~�ӊ��u�����g
�LT^�a	`�%o]�V��������z'��Q��sU	�u��ڹi7���RK;��K��Tk�������ݗu�s>�|o >�5z>�0n]kV�������~"!1�Kʘً[�;��;Fx<���t:��g��`b�{{m_E�i׼��r�O������V雓Rxr�Sٷ!\)���&b�͛�i�;�=ʻ:ќN�����+f��[����3kC��"%B��ZM`�D+m�M\�a���M����`vnk���u���8n�:��K�n}��.�y��kGN�"us�{�nS3Kt�e��\��dKԪ��`h�
��";�k1n:��e�I�ۮI�p=���7�oz	=qu��Ssn��+2Z��'b]�>�|�g$�-�)-�#f��\�(�U�Ų����47XZP������u0ǭF�a����p`��p��]���h"�j�f`���V��t��S�� �7B!��ں�]=nٹ��M����݌��T����탭�<���9Z0Ъń��T�\٦��stܙ�9�p˵����+���(�l��C���*К����{N닇
WS��&��*p��
��f�c8��q2$,6�n2�@���suprH����lWV��ͺ�f�j�;X�=JX�Dj�������� �)��`�]=pc6�(�5�nf�wRfDv�G\��a���]�4rt�;s���mk�:�5��kl�P�#��HL��"-)��@�l֌k�����T]���n�5F[���+������������VQ� ���E>�^�kř6ם%���y5�te2�X�.o�Op�������&�ُ��#Aw*����KΜ!��`N�)N��8�+֗nu^��Z��r�h�|���w"DU��n��xwz��� kG&�g&ߪ��8�۞Gr,����Y���t7G2!O�̘�R�3�9�����=b�r�6NM�����F�ԋ�;Յ���67��o� $��0�7wyw�N�F�Fn��iQ�^�j��6f�,��j��lK�D`vL�{=^�3�Dj�G��
��p��F	�ScF�躭��v����oܑŷk��KJ{�ic>O�Y�%r$�����X<s~�Ǒd�5�bq����j�{n��m��l8���p�KQcC&+]h��(��-�tΗn\<�!��OE���Ʋi'��sf�X���ν����C��p��!��n�8�O'HݼV��f^2��۞����:�6{k��C�8���������U����72�����l�Ne2�/:һJ+���ޣG!T~`(�PZr�1��:���nu_�uY8)(m�nkqf�|�r��hȂ��dM{��캴���:�\V�/Qq��OFk]�n=���2�{w4�!�)��f���ĪY�w=�ts���,OrQsL8�{��b��S0�0��v��+Q�i�M9�M���C�nVMD;�����J��A33c�Izw�A x@�޺o),����x���E9���[Y��ۍ�F�ۄ��IN 3�gu(�����&��m��2T���q�չ"c�[�K}�_/��нzܧ[[�KR�7=M�*�T6�j�K��Ͽ�>~�oү��/���ӭ�!�Lv�{�7�v%4��I���%��������fC\6A�G��ы�7f�Q�Ü�?
\�c��t^Y���A����5F�`MQ�0<�^��o�̚}ս�.��@�#yW35c�s"W_2u0ZE)��p��2f�-��<��a�(� ���vt�ޅڊ�t���7]���E%Q��"�_M>�N�E�1��,���o�y�G�m�b9�]G`(�PZ�ۭ��a����w�9�j$��U��]����h�s�}c���UT����Y[@��n�v�o�&���q
륾X#�Z�=���G���5Z6 �fBl��[���s���#:�M䅸������H��j�`��Ṭ���lWG#sM���v�ވ�5�
g�.�1蜹q|�ص���*P���7PQuo=P*�m���l���հ�2:�Xk�=��8E�ʜ�Hxe�Ԅ殕U�b�������yF*�`�i��F�2JFn�����{:��e����r�q��9aH&TCA���vh�EZ���ɣX��j�ћa߷���k���v�F8Pln���'v:��k���Oa���$i�樚f(L���f�Z�!sҏc'U��m�����K2����i�����M���qaEVo$���v��,�ccH�[h��Xd䯯���
>����KMb��m��9��z=&��x�U���ujqf�����{������v7��a4H� |{�[x�}�-˱���Q����ԣ�9r���V�xj���ɛ�׷��\��Q��5��Z�������v>����s��2q(��Yi%1z�;������a�铹e��{�au˳�[{.�f�7��Ɨf��H�y�aM�*i�;�w+����4x2(��[I�Qy���{��\�'5q���[R���6f7PW�c`^�3��p��خŞx�\������|�w��?.���3�u�i[�N�'D��T�]p��n�?j�.���zۊ�eiN 6�u����_Ժ�<ވ��,縅S4cU��8�x���	7��u�t��W�LSӕ��ճ�yvh�k���pUS�:����^h&�,�z�+��[���%Kǅ^�fcu�g��n#{Ę��-11�s�����dv�~�}0� �O��Z��X6�;����]Nj�	�,4�Y�.҇���]�X��9�(��Rz���wXQٍ֬���ō��m�s&�e���>��z����(C0�� �t�Ժ�M�&DA��:|��L�q����Mb㇒��67']Iy�Լ��7�!�`��\���� �Fm�#	�D�g�m�ᚽ�k����iL&h���l�$�1v��@�V�m�~�������퓆�;D����;���.�m,���p��K,����*0xu[�>{]e��e�{5]�Ҷ��x¸����7';6g�(aGٍΥ�k⃾uuW!���z50$5���~��_9�a��ջN��%CL��ۈD5��î���/l�j8���E:�,�7]O$�k\�f��\<��b�B��0�|�㮨]vp�ZY���bh�5�j��4������)�#	�%X�ݫq�6�ut��4���m �M�	�113x��X��=k`t�;�]׭v���n��?��|�h��[�ޕ٭ŋѱ�1۽�zf�.ġ�; I�׭��a�=��ʶ��OfL��A+Q`��3���n2���Ag���1�7\'��S� �ɛԶ�_�{�/ݖ��č���E�֏�n}U�Ѧ�Z��m}_��ݷ�o@wPQَ��I77�|k)ڰCt2���͙�s�f6"�j͵e�=�u���#�Xͳ9Լ�4&�+9��}������y���hbh���,4e���f!����n�'�ڶ�m��9� {6\^�.�V=��&�1�D1����x�}�GM7=������e'7U�,���ܝbQ����k`�'����B|����߿�>���=��q�h-%/�.�*����;��_\�An�f;�]۽�6s�4mӮ�g�BM�[�3������=��xJ3ǜ�y��s^^�}ޛ�ea��UQ�V�#��n��%n�͍��p�;yk ��.�%��Ɍ���d��z����@����}���"�6MwE�x��}�+cܳT�Ʃ��{p������zh�����:�ڨܜ��e�+%�FRiIj2I�S��E{�|�XE�)�u+.q ��lû��{T �uL�=���]��WʝԣwzT�:�qu���njy`�ݳ7fvF�&� �T��^^*ة��z��7|Ί�Z��y��p�VLj<�t-]�"�	wg��qZ� YM<��%�q	��c��y\`@�:]�dU����S&��zn�;�����À�~���}�q�y��9����oڸQ��Ӫ��鶏c�v��}q ���H�������"�؋�N`��|m�Bm J:?(�i� d~��]�ӎ)�g�h4#��k�`��9��A�������@��K��JE�	�R�m�2"n�34��ٚs�8b��H��bPs�
գ*I�/\6�m��{Jc���$�nXY)�D�^P��^7�S׌%�-|uLx�J�^!���/U����t s�s@��Hu�G[Q����D�54�D2�~2|���kJ�C^D�<{稀7	�牞m�����I\,�(��فL@�����
ŗ b��a�ց+�R[v՛B�� �	"�g�m՗�W�������-k�BY�h�q��jy�t�B��Lя�҉g��G�I:eb}�Q;�C���ܰf��!H8�3�.L+L/B!�hK�-�u.Q�cC��žV�2��)�4F�V��-Œ���w�>���Q�ŖYe6������4�x�0�����e\ޥ���n:���A`����������8x1P]fN���ceh�h���[�����>�{f�SZ�	(m�u���I�AvcsIX �fDAH�hLn�uih����n'u�a8��lN�wt��7�)����4G+n���#VJGf����AWfd�p�δ�G�Ǫvz�ե�~��@��I6�M�M	��MrcM�{�
��3��x����ݷ����?�u#�kp)"Q[/]�Fg�	��P�-Tw ��ۭ����Q��N �JNb�h��n7����	�l���v�x�\��9��c1/�(�ѧC�٘�J>�o</[�x��m8f�]��G�Z�������]3qי��VG��Z������D�v�����3��=tt>��� �D�����-�6��·M���]���N���N)�MI���:h�������uq�Q�����v��:�:��(�p�s�Ks�0+�.������s��d�+���O-u�n�k.ҭ����^�[;��y�L)���"<g.�]�ܩ
��Z趂�N��Ec;�=������]�7X�Z� ������	�E}�������R���&v8��ZJ_rXg.dI�A-������-�G��j31�'<6ێ��0��H���Ao���ک�n7� u��X�0�CLC�n�稝
�7Wf�'m&��(��J�(}O}�7�!q}�����o����KT��n�>�G�Q7&v���&�/u��q�����xD&�0mL�H��}��ί��ּ�C%(i�fkqV����ڶ����F\�]�/5u� C�S��4�a����{���
:� m�K-%��0W=�"�.u��&S �L�{�P�gM���-���O8I��;�{���n�-�� N�#�8��)&<|6ʕ҇���s`ۉ�&%<�r�Vƪ|T	�;�N�k�yJ��/b6 �qN��ڹ�y{�\��@Q�����{�Kf�u(�T�\&�IO{���%�n�,�#��I�Qa��vcq���[�Ϻ������~}}����Z�ܗJ޻v����.5p�&ڭ�T���[�7tU���l�]���*!�/�wx �OY]*�:<{���@&��;�k�bvVQ�a��K �������?	]��1=�mW �3l�z�ݫ���k\wDPI�Ml�=q���*.�]ySH�hlU�nW9�{��Gr��Q�v�N����1�H8�Qa�-�b���f�6e��-���U���+���������J,�iM&QE���9�D���g�;��(�P[r����}�{1��n�l<��6f����qx�E[X y&M�i�)���]갷�>�(�9g��Ȉ.kLv��"C�j��S�LY��{��y�0�7h#��e��Ķ|O�B*4{ـ���E����1laE�r;F�c�{x��\�\P�����:�3��r�C�K�ٮ�z��q�e�=��[n�7R���M�޸�n�k)ƺ���Wwm{
�^��Y/B��[���<�c��F��1)�,�+�7�gb��������
:mf�±�\B�]��b��M_�Zdb�	2��]��6�e��˓N �JNs�浑x�U��x֢L]��	��Sd�7e����}�{����T/q=�l��wTuۭme��ق6f��st��~�(�J:�Ua3���M4�$�on��l��M��L��~��(�z3wٻ���"hu�3br���y�Ǌ�x�]T�-�=v�np�cm-�z�ٗ��N�Ug�|�A8�����8� ��v!U������|z�}g<=]���Ai|����ޱ��]��N^�4_�����A�g�m�X��7l4-Bh�Qܱ��n����e�#o�HE��PT��{��^5׍���4o���(��$:#�"��<v�RBz�����T�to]yk}�P�u����D�o�K'�YLM�4ߟ7����������I1}K�ؙ��������;�%(M��b���^>�C�����C&�A�:�جr�<Ůy\����?��G�:��m���0
�Fk�<�2\v�u�?wи�dN>��������o�5����i�����f[tLnQ�ų5�t�M���T>����fyL]U���ʖK�Y�v��;�����u� }��j7y�i�I����K�ڳiNcq��ms��"���0�3��d�5�툞�M�v̢�a1TToS��K%�Y�0J,2���o}셩����b�V�M4�$������Wf7;���*!�';�ݲ�=t� 5�.#/5@�D��K�G7�a��o�̕�!����4���m�� BH�@��Es_%�	N�Zgi$�A���.�6�C`�6�V�j�MkX�T��qZ�o�-U���kn�V��j�X���m�Ej�*�h�����Z��Fխ^UU��kE�2�ch�cj+EQk|�ۭk��t�J7�\$D|��C Q!�#M6c�\Z֨�X�֦U[QmY��lkV+V6��m�V�Սj�Km��V�Z�UY+Z�V�ڬ�kT�Y���&�cZ�U�+mL�U�j���V��b�EjūU�d�kEj��X�V�.����\TWk�˫��&��J����n��k���۪�H=�?3Ci ��Q��_���u޳����:e�;���J_����'rmh����j2^2�BH���̛���|�`|�I h	 �/�C���a�y�������~($R?���	 G�����N��ހ��� ������G��L�CB�������Gׄ~��?��B�X�u0�@��>+�0Q󌱺��������5��i �$&ВH����5V�[mml[j6�֊���֪+Qmm��m[X��Ѷ����������Z���E[[&�dբ���F�V*�Ũ�4d�V����Uƪ�5Q���@1�����(��4�s�c�C���� ���XI�����>����|�����}a�6Q�� ��H�j������g��a��@� ��������"?��W�Ƣ�g�H��%� ������0}�XO����`�����ھ��|^�ؒ@� �#�O�?����?�~���s����!��� !o�}�I ��?�CD_��_M6�$����?pm����>%� �>��@��RI!$�0eC� �=���@!݄�q���4]�,j�d�$	 l2|�?��|�$	 �>�kG���B?p)հ�o��C6�̈���>��}g�`��>�%�~���a���$�̆����?��I I }��#��~�h�=�>�~XD3i?��R�c����y�}_.�>��?���+�$�$�'�x��(���|y_#a�kg���F��<_Ġ�GO������ BH����0_BHf~;�@I�(�Y�aH�:��>��	��H��1+�w���_��?��������]��B@�;��