BZh91AY&SY�@���߉px�����!���� � �$��                  R�  t       2(     h  �     @                              ��QT({` �Q@�PP  �  �� T�" T�Q@�J�D�P��E�TH���       ��ET�آ��;����w���������G �:{t�L;��<��6�5���҃ �tQ�=��^gݱR���*�D��h�)����_,�S��k�)RU�ݗ��J�o>�y��ڕ����Ixow^Z�=���t�R�/>痢J�e/��:�����k�"R�}$���RR�       ���V��mV����ڔ�e�ϻ�^���4�}w��O��+��;�Ҫ�8 <FxyW��])W���Jy��O�<M)T� z7��R�OwJS��|>��U��l V����J�eP����U<8 z9�T�&�
q4�f��h�������ҳ����Yk��yU/�����<M��|������� Q)�       ���m���� >'��R���y:U<Z^��{Ծ&�|7�<��J����z�R��������s sޯ-P����{�ULM���yj���H�**�N��
�B��/U|�U��sŽT 7��S6�t��G�NX_}���>� =��Ie��A�z=�r�ȇ>���(>R�U       A� ��Ǐ�Y��������@�ɡG� >G���K���e�h.ۘ @рvo���/1�*�B"$  �5O3�1�{�ט�P��wD����4��j�j�����=����e�飋G׸כE���Q�BJ
�V�       �hhVa����Y�{�t�ڧ�;/&(}��j��# ����=��_xƁ���������W��DDR*%J��G�<�|���ϼ��
 l�UX�����_ >�'�[����v8ͣ�s������sx�+��       5ObR�@ �     )�0��J�0 &   00��T��24�� �1��R���H �     $�JBM5R        I�2&*� M#�jz&��i��H��?����~�~��k���q�9U�c�湮~`@	$��?�I% �C�B@	$�����I3����$ $�?�É$���?�	 $�g�q$ $�����'�,����?C���`������������C�ͼ�7�v���p��q��9����-g&ĤM[�Z�ؾZt��q�� �Nsf����Շ /G]67y�v���[��4�Υoe��tT��XЧ=b��6�N�׻9���s����0��ח��l�������ǃ9n�jַ-�ݲ).�Sy����8�1�Ň<�&����mǣ>z�kX#�E��wc�&(�f<�^p����;���ɵ�� ��U����d�\JglȂT.������H�G�G��v\\�K��<"nL$���"e�!�Zr�fFv��v��v�9�
7���횗&�4�6J���O�"	n��޷���e\0�#7��,Ct�z�q��o=���Ӊ��%�&1�=�ش�=�4tQ�Pǽ�`\P�a�*�2z�2r���$q�@+������F����a�8��1���w5��(�v^�v^N	ۯ����v���0f[1s�A��QyX�5e��77m�&Nuy����t@��I�[o7:�w���2��u����҉=��G.Ft=�dR@v�@�I�7k6����}���I ��!ꭳ�M��	l��`G�ni& ��7V+�v����.*��l�=}�.�;Q�p��u��:��/tnl�^W�K9g!����;���Nere>����wi�~��i��ڍJM�;:k���&=S��u ���16�]X3F�z;���+��Om�$�0�:1��:mW
	Mp�ڝe�ю�	�}*Wr�.�N^wX�l�#Z�/����FG.�Q�٫�ǝ���h��S��E�d|
���רl0�)�V�hd�3��(�� )��p	�%�0�N�Dk-�X��)G-��b=�r�Q�_�8�(��Yɍ��2�qG��O ������ZpE贞��
�2��X2���;R���u��Z����cZw���Y��F��"�={��哜�t�F��l�a�����ą���)����l�0#�pROc{��ң�����k�zo}LA�n9��L�q��;�9H$��@�sFV.�5<i���;�Y,Z�a��N(i�5����=�@�eu&��V�k׋�i�~��5W����tB7f�������:��߆h�zQ9�e�Po�� ����gn#����۽��OZՄ���%S��q[�=g �[;{���y��-�X#4]Vb^.��,&d���YqsH�.��:mvZv˳W	b�h�:Ćl��9�]�p�Ĺyf�y:��|,A�ے��
���	��+r��y��ge���:YM�h���n�T���"��N����	ɡnL�׺o��{*L}�qi�^o�Q�F��ps.ٺ3`a���٨<9�;��5�,*�nk�f�$gP�g:�S����L��0J-k-	���3�;��rᨎ�{�%��t�{.U���ӳ]�,j��tsہV��L�Xᝫ�^6r��z���4��y�s���)��;��Ə='��wM��ia�0R4����M�ڔ�7�&ʖ�v���ta��8���#t�ի� �+U�W�I�m�"]	�r.<+��&_%�x_:f��� ���3Wɔ���g-ż�E��r���m�����7�
�.�1��o+ҩW�=�t���ێ�8�0N+�uDgly�f��+<�nf�N�,�J۬ݷ�h��(��'�GpZ(q�b��{�t绳�|��ٮ�r:���_Mɋ�f�=.�D��)��8�Y�J��p��Sz�C���Q����R���R�&���N�u�u��[���Ӂu�����j1Lݻ�i5<9;�����V�K]㥼�����Ӕ�si�����ҳqƍ�̈�k:K����%�����া�r�I�{8N���j���ڶՄv�!C���g��A Lػ)vHno.L��l͜�І��50]�gu��,h⌵t����g��� �Yu'��:�Hjl���h��0��{
m=D9"yT��v�+��ݺ{��i��&v��Ks���M�%�9��l\.������S�к͘��RO̛޽���`�nS�Oc:��Mه�.�H�¼704.���Z�v�|;xT@�NB�׽�� ܃upx�.}d�;`Ǆηp[`�V�n"�Z��w�$�M0^���f��Ts�P؁�e�mͱ�z>�r�ˉ����2�׍�]��,��5�(
Zbnt����y���[�0oI.�4qf���.�o� sі̴U�6]�D��f��m�VZ�.�Џ=p�]E!:��B�P�ٗ�ܫ�׏�N�3ל�8��2���5��	:j=�S#��)6��ٛ������0�\�q�p�3��s�/��h�f���LB�|Y9sd݂�Ý&4*�K2��\���Σ�#5�O+�]��ls���|@=ڱnsN,>�.�Í��k�2:����)E�����e��ܓ;�8���dhL�䭦@�eo��'X��n�s�s:^��EF��V,�I�dg���ئ	� �Jb�2T���	C��=��C7�;5���v��J�yf��n,��~�]��Q��=�.����9b��w��s��,ւ�E�6��HPv!�o�rd�Z}�g=�]�FܯlCu�*ZLۜ	؊oF�j��3�[��hn兡V���z�N���#�����N��rn�Y-��ZMK�[xQF�ٸ��vX�-t@o�b�Xtl�Ӝ��*"\��VFM�Nh�Ƙy���<��iG�;A�N��I��@O� +�G7N���sq������jvou\WSɊt-��C�L}7|����jf�Q��;�Gf���
���;d=zw�ye�����V��{��V���F�F]ZE�T�-�@�rW�s����M藃��i�F�A�f�v>يd*H���A����o9���8t�Lq�L%���t���ݬ��7B1��D�iB頖���$�cl=�E�
4�\�#���iޫ�w����(�!��r��[�2����<��ʦNSbf��i��C�<W���5C���z��q��-��D�du{��X�1�FS�\y�Lk���*@��,����2���k��w] �![b��\+z,�ˤ�<;�
;gq�9j:>'.���/-EghD>�.k�r.ΈN��Oz����-!F�:9BS�㽜XC�G���ovAë�RӸ��00"�\Ľ��)ȃ1�5�}]��Ԙ��o�A[�xeއ�]}�Z�!�jI%`��k���:.9٭e�秀.K�Y)�y�eQ�U �Z�D�ᓒ�,�j�M�q�q�9���e�Cjnc�K�j
f�[�h��&�]_|B<��2R�t�Fv�\ѮW���|F8��µ�wv].72Atq!�/�iTK��D�;N� 캝1.a/��;w`�`a�F�v���>���ǂ�uz��bL����/m��54� ��/���f� =.��`��g=��o7;vUEt<!�h'L�JQ툹d���%@��V�kp<=9#�m*�%�+���;$��vs��O.<�k�f�\t��m�
5-}�GT;a�k7s�!�&��4m"	���^�0i|�s]��Wv:{�OK�]��5cYkݜrp{��j�7|%3{��v�G�w4�l�ڻ_C��>�F��Q9a���.�T�G��@��x�5�ƴ�#KG��U�t�LΤ��˻7���H�6΃f�ذ�e�(�g6��7�g��&Iچ�hᛝ�4���"w5�wH��3zv����t,�u�ouÎsOU�H����{aw��8�pwDnt�����U��6f�z��L��Gw���,��T�Β�v�w���f7�v<]w2oA�b�{Ô*C�-�+ v�&U�r�dx��^;6�Ȯ܎E���hK
5'��^XX2�A,����2ݸ�p���e�o`�w�zށ�G����˱�Bl�������k��ђ��s�1̯G����rw5bW8�خO&��7u���je���YX]�0oA�J��[ٗ����{f���Fmj��B����8��s6l{F���u.K��Z�ưMM �q�q�"u�F��d��v�AT��6	�9�M��v[�V�C��f��B�}Uȓ�cfΉ�O�/�K˅K|OoUN��J�477{��!B����Nͩ]�n���v^`/n^q��|o7-(�ћ��=�)�q'�s�<0Uw���3���ݴ>���������3��+��N=�riJTf�:Q'���[���1H�]]{D/Q�0p�|�T��1�.L5�'D�W�.=�z���l��jcB#�?�lv�� ��[��� JN���9BC���3����h����7�C���=Ȼ9s�ؚD��0ZŦ�����Ȭ��NiW8'U���.�����g� s��ϻH/�vҞ�miq����Yڊ��s��}���3��a�5=��a��`����Ihv���j �����"QZ͵�yƴ3��G"�������WIk�hU�Jo!4��w"����>���i�/�p1��t��í2���m4P��1��qoZk��x-��F4ɦ��ܙ�җ�,1Z�u�k��w��Ur�[��:�Օ��.Ý�s�	y;8�����ҥ콵��ò�Xyn��{!�.!���>��:� �a� ���8`�9�=]�K��ź��(A��s�w6��{�ܠ�������W7e�,����سdpyq1���u+u\c�ң/���W���\�Z��c�R��Ȏ���w#GY���f�.�D{��o���5T�ה7ۋY��9ˀ���	�q�!�똹�%�w����nn��g���um�N�L��V�gNl�Sx>��JO�>�aÏx��,-;�8:�k��nm�fM<Vq�N>L� l�����6Y���q,�޵���k�L���'�N����]�].-��17~ch��,Z94Vh�c{�a@�sN�k����錞'q�&h͝�A�s�'+�����I�qns{����>��Sb��;�!N	�٫�`q��*q.�-�r��&4�E.�;{p���@��JNp��gQ8eu�}�c��=��*��*s3V�|�="�Ct����4mN-�pD��MC��q[���.�eՆ �T���t�.�����~�L�ռ	v�&��ˊ٫<sr�YS-�p<y�0��9�����/^�������Y�j`���,�����o]��͝���*�Am�ph��֔�K��d!W�MP��Wkvq�y��+yn�ot�,�^&�	N%Ï��U���������w�rNQ�[���M-A#�n=��q��@΀*��4�T����O45�;q2_b�ҭ[; 0����#��\V��7�,��+u �n���a�����X8F,�6oS�oG�r�z�E��]RYn�7��*��|)�3�
�$$ͫ{�mocs7��2f����
e�Ӑs���ʮ-ݻh����7�u�R�����@:�q�L����YFh&���g�
J������V��*̓sdM���!ؓ:���ͺE�wA3��}��S�\Yq8��ݵݘ��n.��Wp˽{n���ݣY��9�Ú��/4wY�vx3��u���pd^���Fu0��;�5ܽ���%�
�d�o	2�g�9��Of�ZB��	o�#��9�kz<��y���,��G@�J�{(��(��z��V2�h�i8`����{64їSo�K�u(�>X�:��sZ���n�k�7XqŃ&;�e������ø`��E��R3[W�*���t;+9�LzX���1�j�ǎqw����ր�3B�)pb<��OY���Z�Հ�7k��䷅����h�R9PN.]D��J�)�T�\4]:�ǵ�n�Rtۣy��I'�Ld�^ω�C�Bd�:��o>��7�S�s��=�=����N�^:BZ��2ϴ��T�w"6��u�{��:�S�L�v���-y>o��:@K�\>�㋕�����i6��kl�H�6[��o&Ňuֺ�{�8:��t�}W���-B@vQ��l_Z�Fn>K��T���^w-���2[�g!��Π��Qv��p���}�ִ�k�l��d�z^]�pJ�KZsp5�y,᳢٣';wW+�q.׫:��J�ǮR�6�:�>�<����Ţۜ�J�������L��k�[�7���B�-���t+��.�yw1'i2g3b�Q���X��`�c~(ۼy���z��"�'.H�Zu�ya���wv��2��Z\��r<yZZ;��ʷeڜ�:gi�ɹ�k��\��O}&r�C�}UȐ
�Q�`i}�p�-��E���r��ۜ�U�ZDͻ�WtZ��X4r]x҄�Xn."�R�[�SYy��������&����n�pܣ���N'-�rˇCe7�(9�ģ����Q�� !��T]躬xE��W$�;5��sU�Μx���#���J�>�і�Qډ@JCCr��<X�}-Wj��x��!�w,�S�˟tKW(2
����k�&�FW8�@w���I�}�^7���,,��n*��7E�nt�6+y���w���^��GӔX��b,�Q�g;�3��}��u֐g���\�D�ٲ����˹3k��jÂn�Ȅwe�����7���[&�j��R#O��ۺ��#~ۻ����p�(�T�ⱐ���X�g�s��ߎ�}������!��؈&	I�)A�l�9���\cp7���uk��n9K����c1�9�<f����Z��uɱ�����|�������&'���돰�{�ʜ2n�c,Ȗ5gv�'%g�iwfx�,\�<�]�f�{{N�]������r\�\v�X���8΋��.�;ɥ�.�o&���=Y;n]"��j�t�o.���m7�uVG[>���z�\���:�]��+c]Z]�g��^�؁��v^}v�n:,���ч�r3q�-�'-��r�e�����N�aٗQ>��5bv�������s�&��=�r���ƈ�d��:� ��l��;�:��� 1��wv��K���qN�6�;=�5=s/5�;Ϸ(7iq���N�n#q]sl9z�Hו�L����$��]�����NlM�G�n��l�^[k����]�������`uA9��m�`��7�I�G]��4@s�O\��u�tW[�/��S}��aqG=tqA���n�MI��.�N��e�j��{%��y(앺�s��r��[����X5�&�]�g���N1�9�ڈq�eՎ�2������������Q���k�P�^��e�q99��mm.���'�E�����9n,�����Ѽ[	�ܼ��3��u�p=���T���Ł�p�8���b�*]�<��.��u�$��h�v�4�[Ǟ������ob�o[q��f� hV�x��j3���e���;��6j�Og+� _װO�������{Z.����jCc6y�$mnq��1�6\[D79۞[dP;u������`�gg��l�i�nx�g6��\����6�y�1��un��-�7;m��!{]bᷦ��n��d�nŲ	m��0"��`�B>6�Ѭ�9|;F��_RC����m��'%���z9�ӷ7"��r�g\�-�wK��Յ;G;���D�e�<8�;%�^	���G\��9�W<Y����;v"ã���ka\g�l����ѨH�<;�C9�r;^��݇[v�v���d����m�1�����ۨ�oIļv�"�:8���9�cYv�܇�u�7\R]���ͻnG�����s�l�K/<��᭎��<\Oh�9�v�v��93nҶ8��q>�F�t�v��m��Zu�q�hǟQ+\6��Fn�g��x�g<h�-��j2tʼ�;��<mjRq��q�dXu��[D�lZZG^�ա����]p��e���Om�n�f��)��s6��������~Fgm�<a���n�-�k�x��fݝ��of�A��g��.ѼL���%o\��^��g��l8��~e;_g�OG�/V���͎�.qY��E:������xr[�X�:�9����y�5nM����3��I��Mō�ݬ�c"�Z穮���:떞���3�g���z�qY�y�v��nB���v��5�E�{np�<1�q��O<�:�wl�Gu�s�Q��x����ɮާ��wV6T=ڬZg����՞{h�b���m�������8�5�p�����X��7tp�:�9�˱&�4#�Ԗ&�6|��{=Ov���GWnz�g��ϧm[�ۜ;ũ����Iڟf۝�G��X'�,�4�v�`��xE�b���*�;aQ��ƴ�8{���=�u�����۞Y�na��snm��j���|�϶un�C�����=��%a���[Sу�[v��{k%sڌ��y��L��N���]�9M�ζv}YK���1�����|����ux3��ն����a��<�x�������3���q�ܯf�޲瑞��\���:x���8��6��5g��x������x���ۚ�n�X׶�;k��q���n{CҼ���ݻ#�Әi�������+m.����"�Su�pv.�g���\��!�g46���۳�'�hۮL��(�'��=��0�n:��v���A���μ�L�6�!a�J6��r:.�db������!vζ��@wd�zv����=�<���{<Y�nmmϹⱘ�a�طS�z��#�X����&Ѹ��B��Į�7V]��$C��[���a�/=.�h*��q�X��q̓��t�A�i�ku�Y�ŭ�o#�L�X�>w;`2;�A�E��t�g\-�[��Ւ�r;ƍ]ۻ<���xF�v�q8v�\���C&���=�u`�yt�����/t�7���dwenw ���@���6�*9��oN�ǎ<��c\ ����^�,��è�îL�����R�A�Fv��k0����v��D�3�`��õ���9ik�7����K��wcy��+3q��U���˹���#�WJ�p\�
=q�u�rlH�z;�ny���p�>Ӂ3���c��^�Blji܈�b=Y|����r��Q:�6�c��� �gZ�3��zF����j�vS8�;;���6���q�#�쑫d����}fܺ��k�F6cq�nq� ��ͳzy�;0��0��c�ֳ,\���v�� !WgC;��ɩ�Wc�n�����ˋk����1�/Ork�y�ց6�<�M��=��չ�s�!��:mXә��C�u��^{'�ڮ�k��u�õ���ۛ= �=v���.��gn��<��^�p[�����s�hM�!��{��pqG3CA��� ����i�¦�m��竖ݳ����˷�aEn�v�tm^��F���������Q�W`���[p|���ˢ��uɍ��kӵ�Se.C�ޫh�n���W�t�Ntf��B�ѓ�.��y������^� �童{-9���W&#-�K�F�v�m�L\&��W���2]��;X��m�ݾ{E�3��e�����_��7�$Y{]�796m�m��9㹼�'F�K��LC̩��ݐ��s�oGl�C�� �φw\u���Wi�h}i
�Z�,����Mi��D��62N�_=Ν��S;<ɧ�����n��[^{�K9��ls�Ǣ`I�ǣ0����m�
b��W�LQvN�Q�9tp��p�J��h�ֆ�].�s����!�WC����n�ޞܼ⛍�:��VG��r���=�Xm��xq);tF�[���ɭ�9�p����s�v��k�WV�a�;73�C��]�\�0��׌Nm��9���ѹ{U�D��On��A��]����Nk�[Gۭo�\�>C�sѸs7]b]	�\�i�#�]��K@A�L�8�g���:��̹��g�Y�t���n=�a^8t��-�7H�q�������+�v�X�L�W�uێw�m�\�w+�,�m۪�Y�A��S���<�<Ϋgi�p
m�C��6S����=�㳲�kǲ��I�6�ڎ7��� V7�k�3�-n<��<���x�0h����Q�wW6�K������3u���m����'6�Ǣ��u!�+���B��f��ܖ�v��iݫۓ����Ŵ=��4n����nv�����۪�4�(���r�X݃�r����s)����\m��[q��a��^���v�n9B#M�?|�.G�c���v�=��l X1�n�7�d	v��',�ݰ]�n�=�.��x�lutz�v�1�ƣ��j�юL�����vc�C�l�e�t�g\�=n��l�E��qV�4r��.���=Y{�˱;�gk�n�1����z"�5Iݚ��:6������y�=���m��ν^z��;��[X��㎠K�!��m���<n����c3�[+�[���W5�-�]���C��Z�Kh����(c75�n����]�8{a�d�n��yG�s������GK�����k���/9�p'c���xeҝ���a��G��s��A��B-�<���9�㹒:vg�uЫ;s��{i཮���Y�9�ӗ���m��j�y�x�䂹�.�L��oNw�x������]���ֺ7l1��u��B��ݷ���6�κ��^,��ͦmJC����\Q��Z�HO�|f��Q�0X��7�
8�]�ƊwC�9����̈́��;ؓ]V�7��=	�]�]�J`:����a��B�۵�������;��<���[nzH�Zn�5;JmO�N�I�/cű�ۥ�����z���_=WKmR���p�.dB��\nj2�V�۷1[�^/b=�W��&xn��� �u�޷:�ʼ��K=\��T�WvZ��c�zwg����#�(�q�<�5OZڣB����m}]��rTlv���Sq'[mǜ��kxm��w���{�M�v���(���k������,�s�s�g��Zn4m�����8�jt�Wk=op�V��b�c��	��8C��c�1���ێ�V뀃V�݌��"�s�W��9��v1lv�ʵѣ���\����u���U܏��#�N�m��鸻�n�q$�v���]!�::�[v䌍v������֭��nqv�
���ۙˑ�v���\v`��װu����pN��v�}v8�6�<;ܼ�[y���v�<����9ƛ����{�Fc�í�l�gI��9#�nn�ع�.���t3����\<��{]��x(�R�k���O\���o9�-���ۭ�rb�ܯ�(�8wc
Ɯ�#p���y7�;�y6Ħ�%�;�w}������DwjP^W6��\�Jt�r._m��1��{X!)��`�mv���;��LU�v�d��W6ugW�}�>�f0o�6v��]짞��Ί�Fx��6��Li��$w]9�tt��(}���ݹ��'9�有�׃����.��ۆ��=����I� P8�{$�Or^���A��A�`ic۔��R�N1����l{	��2:�z�k�vCd��v�lok]�v��svx��n�C���[��|�\�Prm=���r��Drj+���n��s�i�|K�3d�6�X�C��췌u�ds�u�e�����Fh�RF�2ع��S�=G�7o��C��;q�Σn���Q�oN�5�n���6�q����L�����ƻ �h4r�m����y�j��z[k���8F���Xa8h�u���V���DaL ����F�.0�xZLXɞ�x�8�D���\�:0�b0����]t�6��ɳ'1�`պ�>�q ƻ�� ��Ꝅ��N8�硨��on�<u��6�Pbh�.i��=«k�hwI���m�ؘ�b���q3_� �I�0$��>����#���W��S��L���3k&j�d��ű�Sڌ�K�7����?xRD4�����2"խ����-�:P�ڸUf��`�h�5�M���F���(�l��F���#a���"B�z'L�ޏ��y��=�U���Oß�����]�G�p���<|������{���l����>ŵ��E۴/{/��3�Ti��%i!�V8�N��&�ѿ������k�R�/3���Nf���	;�*��Z�B�5yC�C�H�n'��y������u��w�R�27Uni�]�o�ۜ=v����Y�e�_����!����
�c�IB}���^���6w�I/w�a;���y?�����# 9{�|;nqY|�{B-B��c��|ʶ޾�+4B�kɀ=�x��}����qM��j#�ōzQ�ID�֬��<�xp���y*�>���`h���O6>U��5sd�k6�����Qn�2b�\��t��7��T��STY�v�U��J}�U�{z���Ԛ�����Y׶��p���Q�_l3��N�Wf��qzhڼ����s�PrkԻw���������z�z�r��p0
y�%�GR���3��g����VU}m�<:g	�:����w@6��~���r��?�����.�@t�n��}6v��x�b��NKK�Ͷ��ߴhwV"^N��Qt��' �`�v��{Z�2�#�3Y����6���?+�Z�ҕ'1��]�N�2�^�'\S�ɭ�#JAf�Ŗ���t�m�
��S]ΑG(���-/��D�������w 7
�@������M�n�%��]٣پ��Bw����t~Hb�5�����bt��1 ^����>��G�OD�4���;m�~�ޮ�\��i�Wj�GQL��9�����ۮ�D�t���7�o:aݾ�ڜ�OlhjȽ�pj�&�C$��x��R���ozz`�����a�h^�W�+lKX��+�,�a:�zϯ\y>�=7
�y�m>��{���=�z�]�F�C����N���q����w��������K�+�$��V��jX��1�N���>�����7ۂ������k�{U�����.��D�b_��eO
���gv��ݲn��/�Y��ۊ��'$�{SVm	c"��f����n���^�h�hb�ͭ����ˤV�������޸	>�G��2���F��sgeY�EuH�Y�s�o��a+@��nvR�@�ū����8�ǹ��_5�5
��h����`ʡ7kkIĤҶ�b���U��.]����I�q#.�/x1t{-���e�������~k��+�<r܌Z.��|������Z���Tn�����y�+�������כS�݁4�p��c�p�4W|9�&��ٽ�u�/{�"h���9��6��*SJ/i�]i��C�KZ��;z�6`��F,Au���sIª�rn�~�Y�Z�`n�W��{sp����AYu97'��|��^��N�pf��$��^s���g�{��`����ٻ��РwUǋkswu[ĠLJ��LC�3�9�WY����Gœn��R�q���a:f>��Č����o��D_���{=���{��wtc�<����(�:�چ��&���ѾO������ބLv3����bĞW�o��e�]N������;��*íХ���������;&A}2��P˙",�{-�"E�E<8"�3�v��䳀{���!a��~xp�����D���n�so86,���Q�g.�h?x7�}r7�#�Ӈ����k��ّ�����8�TR�� ��eBOm.�;��ϻ~�)بF��7��y��4+�h,��f������t�p����f�U��Z��yL�f��Z�΍�]^�b�q�G7�Žz����m�y�U�w����sN��&H�V�������O��w�����3/��r�7'��u����|����b�6S�{d���}PQ�f���S�����X{7ٸm��V�ga�V��:�|7'�zh����V������T012�Hz�����v��8�~���܃�G�j[5�{3��[%�8�Vƾ�!��Wy������>��SO{C�3�`bg���_`���m\���c4Tm#v���:l�#�ݓ�'N���{KI�H�����p7�i�������@66�}h�^�>�s�E���k�t5��O�3'��'���}�@���[4��N�>�O��7�DavB ͂��q!5Y�p/ٽ��z�=1����'o�^��,"��k��yq�C>�륿���40U�*Y3U;�:``jL��/;[�z�y�ۋ6���1o4�P�Um}q����z{ۆw�����QA�l��[:ƣ��D�&�%�==��{��}�H��I�E�����N:;�֬ރ��(��>ho�����f{�}��G�A�ܫ��������!b�����{\�r����Q�(~�ݝ67��ls����fl�Z���6��<{H���y��y�UG����jy�yT�
��_zd�}�(����hV���ٵ.�@w��v��_���
��4�)��u�!{��l��;iZr
�������׈�KH�тI���d�S����:��'"��9��.˽�޳���/���]���F
��BJ���&%m�ogw��R��)�eΐ�<���J:v{|�П���G���-�:eö�$:���=���J{ĭ׎��?nhO5��v�^��o����w>���9�F7.ﳐ}�Y}x�B����b`�U7�ڸ��X�g�9����1�}3�MY�y�������Y�Y��2M&��m�E��S��n�rs�	O��;'���tGx�O;��9��cO�_���̼���F���a�Q��V���3��Drϯ����j<��s�v�|ǗxfƉ���XB�'FF5)H{j�!�A����0o%a��"M��U �Xʙ>�}a+O^��pǰ�N==�s������˜nښ�R�|��`�RQ|vۣ{���O3��������Y�J;��c��B��Ӑ�rs#fo�h�.g�]�^nH��U��*�`�S'�=��tC�B5��Z�^��ms��ܨ����:����&6�u�C�^���=��݌�Y�*Mz3�p�G�z��焸��F����l�}�2������&��c-Q;Gܯ_�]�5�Ga������H��;��`�6�v.a�VP��K���{ӷ������[����i���ew#�3��h�"����Q��qot�O���)��s�g�ޒMGXՔH��Y��c��i\TUE��a�Wc��n�rn1�8h�x �M5�[v�Aj�dY� �w0HA%ޱH��Ű�=!��;����&���n[N�Lv�i���T+�}]���oD.�����Xq����~9�6��=�[�q��.����C�1�ꂯ��qly)�����p	8�nFވv䉐�wllm֤��<�ͦ��~S����N>����;t�l阎v-��g>�������疄�� �3`9wj�k��N3kF�R�̡�+R��N�-�j7ca���"eӨ;�!b�Iȋ�
�Nf�a`ǗW�<J#M���P��9�p�=���;/-0d���ĸ�=�;�G�?c�8^ئj�>r� ������c�3�w�]7[��۸�>W�W�z��#)3����g�����&�F4��x�6�ĝP�rc(����;`���y�=�K�[̫9/�ͧO��c�q�D�w�v�~�.b��>i�om����%ɓ�[x�;�B���4�w�L>|��9��D�������vC�jy�P)d�B������"�^늱n�>�Iܰo��w�C�Tm� ����~����޾f�}$Z��1X�ָqᒜ	g;�#�1�a���}����헜����N}�i��l�w�N��~���;p�c����-��\	e����pE��x����=�]��zM���<���:s��=6�{�yz$%����7<2n{�i�2���;]�%2YR�?���my=��W���{̟/7����k�������@����r��Ũ����{�k[�3f�^�F�)������w6������ӠSB޹0����0	�,$�Ҍ��R�.m�6�N����HCF�x�	C�o��U�V��d'��h�F���xpW�$���7�rj��޼=��O�[��S��p�D�x�|�3��V�uk��[Y�"v1jo���$.f��$��>ȩ.Ps�	�\��/P��C��f��z�]�l�l� �nx̾��_g�#�t�}w�aF��F�@�U�sIы&�	'��qp�t���zb�aw����� Iz��ڏ�h���,���3��`���U�󦩰s�ޖ�0<�o�ea�7d<z��8�i��;��i���/��]�e�� �[�2�;o-�;�N����yhC<�ξ�8Q����]���c��L	�t{�=��}��,=�N1�.X1�.�P/5��Eҫ>^;���}<O��w��=�n޾���רU����������F�f��Z���C���O=ע�ɹ��x�(^'�!Trܾ~���o|�%� �9�A��e��g�{�$�#���>C�_o�Ϛ��y��r�T;���n�9��S�<�QV����>�2���|�$����1ѱ��U���e��Z	�RW�9��h��Ɵ|���N���e��[�����w�95��n�l+��Ñܟ�2����:<1{�z�MC���x���X�����"V`i;�[&���'p��\;=�N�nM��:�|�M���Nx�tOV%��	�ݦ%\��8;��wh�2?M,Du�H�Q��?C66ؐ�fl4�#�j��cu{!�� ���z������;��F����g7�ٮ�G���K�j��(jӱ��cQ�J�ܫͣt��[��a�~��;�� �bz��c�jo����.C�͇-��<Y��v��l��F�rٌ�$b�p/qF��=�[��^�Z3��%��7�n ��N��L�dJ�.P����7M8�3�'V����9�_yw�P�{,*�Y����:��Xv�Ǖ���]�kj���P^H)���n�Ég���}RR` sի�����B������;٪�R��ZR�f� ?%�J��Wڲ�~=zeW��\z���%��we;�E����B��Y��ÚhO�_�ʘ?b'�; !w7�-����i'	����|�8[�{��T��̎��h-�������3�w���'/�g��=|3^�.{��>s��
�i�⍍T�Ԣ܃Yw���!�eF�;�s{3	�XI��a_ۃwT۝��;g�}Z��Fs�{�lw�Vȷۤ8V��_�� �����s}���6�"�je�����I Ưb���2�>�ɾ��O����D������ԟg��^}��V,�<�n8����2���_�/w.}�N'����������M�=���7S}_"�隧8e�t�6K[nTm�w�<+�o��x6t*��zjg(dhJ��cnf�����*�I���������p�*F����[�lg���V�bX~�֟����e�n�T��M��z�����ᅮǹ�q3p9iԍtn�*g���1j	�_7�'�^�K|���>��✈�>�>�e�<����N#�7��gQ*��?P�&�n_nj~�{��T(������V<o�d/�}�{�v����/v������?�$��>X��۽�����j�\�z�Qԧ(h��-�wF7Q����Q�~��v�qv��n�=�Tߟv;��8��/?g�ӳz�+�1���Ѧ&8zL<@��"�u!mۉ����
�L4���{z�_	/d� ';��ml��ui?���w	�}��71���&��9�-G�T��f��tpD����W:�˫{{�̷�me��;���Ǳ�خ��h[�8z�^�,��i�C�r}��w X&�5eY��B�x��p���ݗ���ݓhG���Eضli�36��Pu))��Z�e��H�Z�L��ޞ+�Ĥ�{�~#[�/�?!k�{T"a?h {��'�m���7ǰK���Ӛl[�\�y٪BE\�"���P�n�_{���=���_VJV�@����g%���͙�1r�'�/,9�b|��0ܶ�C�q�.�(���f��j��6U�թ���`&��A��ΜWxA�ݝ�{	��KX؁+<�Ḥq��Z����V).�s�^�d2���+�f�s�#5����SOd;�*�2���Sʁ�'_b��Tf��G{�'7���ߏ��M;��Z�(5��w�������sB�Y0j:Z�&y����C�.�̻�Jtm��=��/�<�o�'=5�b9
s���%oq�ӶX�+5�tJ�l�¦	"�� a��Oc6���:�B0��/o,�e���љ�&<���G����Y� n�$^Zݞv��l��|��8���>Y� �}p��Y�7w�,!�}�������e9��U�������:�'nx�W�a�{
s��s{tN��ӝ�@C���G��O���^��=E-��&��C�i���k2�NU��1���!������NJ�����<�-� {��r�nZ{���5`�� ֶ�N%^��>^��޺�Y�/mn{���� ���ަ�s��V%��������vIE�۳����� ���n�U�|�\��F�Bv��1�"F�r4K��,F���7:����3{��b礛�`�@�j�������xl59u��Ͷ򛲃ۋ˟���~���/����g�9���F�`͞���W�j��ݾ�&�N�GӰWV�;�\�����3�UzF:C�ӵb!{C�J���=tz{y�#p~�<�{W�2#��qgT{��J�c���9]�5e����}�x�����cc�v"i�$���77
��N��g&�v`"�)Sp���_F�UD��K.��+>GD�M����B�=_{�_S	y^ ;�=��ăܩ-�}uE8�?1�Z��_jӞ��ޤ�����x�Ow{�.>(����"C.S��HNV�]eT��m%g0kûIУ;�&~����g�Z����O� I$�l��?����~����~Rk򤤥
bR�H�����HTVn���W.;u��ro$G��=]��
ʻ��Ng�&zzo\��Ů�T�=��+�]�/�{��y<qoc��v���s�7y�q����Aۜ���`�zyz�d���m�1Vn�F�7�wǳm�r��n�6F�_,�����^n�.AN�gg������G��Ѻ��utlb�`Gi8��1`��ے0�g\Yc]� ��ϵ�n.1i�+�۶�n�v^޷V���b�zq.���p�89w�VN-s�/oN��4vp�gFy���k�]���7lض:�f��6��cki�yݮ:��]���y.ֶ�N.�9�NyV���8:�Ú�ݱ�c��˴�O�E�;e��:�s����gm�JlR8�q�Z�8z8<;�`��rط;k��x魼��9��vG�������\dxⴣNŒə챺7:�l��� xxC�3TЁ�A�E�e�k����\7�P"�s�W��U�:-�w6;\.#���n��ݻ"�n6vҜ[Z{yu��Е+��^��/6�/;z{t9W��۫���բ.:4��cb1�e���v��[�����.ީ��*oj�v'�Ƴ�xp�ƹ���������>�[��9�l�����ob��*N���.@&�xF����Q���R�㓵Ǟ�m��7[�N��ڻ)�cMǫ�!����f�5M۰���v۲w$\�=Y� ܗM�ų$��L��]��[��$�v��	x���݅�M�y��g6�׺��N�x�ܹ��@,�ݺ�n�v�t�D�>z;x���M����tY�j��9���$�B��h�{v�c�{l���Ge8M ���ĺ�v�#g�xhvn.�n�t=����P�S���s�Պ�l�w=�j�r>�.l��wk�>�۴[��;�S<&��=��ls��֓��ֺ�`#X�j�z�cO�vܦ����[l�R��t��r�������a��|���l�˞�.�n&��˵�7s�	r�\����/��W��q���~nqf�^Y!�c|q�`R�����y�,-���OK���X��B=k�^僸j�A8�Kj�e���ݺ�
�L?�҈���|s�r<����b=ѝ�{\����O,N�骼�00o�5�}x��o`o������gVZ:�:8R�	/\ۻx���S�^�8��Q���Haa,wFo��c7��
�}s�@N�J%
����`���e-`إBS��}�9X�4�G�t��Fx���|8�;|4u�Op43`��6����ތ).�Z�R���i�aC�����ݠ`�d�c��"?��1�������ǗF�S�վ��wr��Oۨ1��Tʐs����q2��wP�� HJ����7s�`ȃ�w���V/�łAXޔj��FϝB��`y�h|���f���8�A�M�y�鸧݄%�2m<�sq���>@���{��:�.H,'�jBX)����)�@כ٭=��kz`�W�u��P'� �c�p+���ɿ'ۺ�#��`#��IX'�N��J��'d/�j_�+_0�(ڳ��&s
�� ��k����#���2C�o=0��&�rgMH��@`Ÿu�ˊ�� ��I����b��iBف��+ r@��.��V�z1 �OX�J��Fc$%��n%k���B�	�2�[���R	3�1g��={l�����O��Q��&0�N���U���Q�i��+z+;sΌ�v��x�v������:�m�i��8�7�٧�g��z�t��R�.��8*�<rv�����{B�D��F��GY5v�'�h�݊�O=����[:���Η��̶H��ڮ���0sn��n������T�����Q�s�o,q�wO(nv۞�X8n�Gs��vF��j'!��؍��H M")"��N릌�r�w^���~���dC����7#�w(���*�a�&��9G�p�(��tit`"��3�=����E��uz��6��#d3�/�a�#)BD�)M8w�
� ^K�K�R�k�F����>��5!�"n5���r�d���p�]�� �Y��wWp���)PnD�ɧ\>g6xf+H�Z�WT�~rw������	�[�P�+8$J�}����B̬kT�&�7x��w��|�p"B6Yl(K��袼s�������������p��K��^�rU���#����0�ѕ��wv�ԓ��^���d�i�"T�Ɏ#�e�$�ڇ6�]յ�V�X�d�wOJ�[�zvg�����ܮp7��S�4�����*o��qw�1Z��2&�Q��x"�j�u�ƛ��<-V�VT����Ό��uX�h����ϻ�}
#���,��� ����	�R)wvh�{�?��w3����P�]����i8�FCM��^7�z:-ݼZ(R� ��ޅ�V���52Mc_���f�M{���w>&�K�[wn�d�$�k�L㮎�woWT��d#��
iF�y�>/w6tUS]ݷ��]���A��}��%�n�	 �!��j�D-��*6����e	ѧnε���[��v+�m�
���̋��xv��W6�)��v�mDp�wsw�]ս��0Rh��p�L4�pi�w�E�|>2elr�T�]۾��\�� }W3��P�$�m�H�qn�꞊UNf»�9��\�eG:���n�>��7�.�L�K9^
�n��h��p�HB�W�'m�X*�T'9�S�[yKoT�^+���>h����F�QT�"J%Gvỻ@���'�)���D���nڇ��vp#3 �J0�)��9ϳ1ێ��M7��?�����gN����E�f LfAH�
��{F�7�}��j���S޿�vl�P�e���p�����J4�/:��t�[�u�c�Z/-�w>�X\�ct���u�^��2!eDCF&�m��w�ӳvq��J�üһ�>̼�/�Ӧ�z�JTY�jpPv��Y�W���v��L�J���9��'2bu�ĴXjB	��4���Wuo�4�����v��Y�x�!���l1!�6�svoj��w3����~�V���6G��7��C��y;f����}�H8쌜�"�᷺�B�wT��;J�]��˨����Ʒ�I��;��9�~"�so���z�QQAH��\!�4�* �I$AR$�Z�x�w6:���h��p�$�i�x�U*���%�f�����n6gRU4�}�ӨP!*a<�@���q�D��W���RU���v�#��)8���R�Q��û���W���tR�p�4������ss:�U*�qH�eȉP��-���w����W�=��J���;�S�8"� ��Tq.!(�!�M�wV֣�i�x�U. lf}�&�M�"�}���G�y RRCJ,��M%S\ 8�`Z�x�DR�p�4����z�Y�M��G�j)�8L���sMQ�}���fN8�IT�v�M�L}ʋ�W?~Fs������N�;�*�N�FE�Vntt�E>8���1���A�wF��ĵ'2l�r9��]kKY���/�ߒM��"���846tѱ���8��[s۱�.h�Y�]=��kp�g��pn��[�bn��㱃�o\����gkj�bz�F�.L�c���h�����s�j
������f�w^9�c>��a�n�M��ٹzN:������?P�kz��{Y�|k�óƊ����K�۷]k���\�5�lӘe�+�㩻-�fk���Ͷ�{�=��`��M�ۜ&1on�ۻv���J���'f�.�{r�WO��|n�v�{�2��5���z�����8Cp�E�*(E)�w���k�4�Z+�}n�Z�*�,}�bp[a@A��V�^%��ϥo�xd�k�	� �4����'k�L� ��0�
-�tޮJ��xU߇�<w�2m�OU4�͓L��M�"��j�N���.�:��Z�����v4�J�����Z%T�Y��wk� �&�%kv:-ݼS�)U>��@����m���vF�]�'qh���v���YV:7\p��C�A#1���q2�dDR�Nsg/�ڸ�M��n�{��Z��;�.��𬌜HjCI@f���%G��x\�"A'2�:˕�rf �{�+xD�)<��"�d╺P��<�^�u�p�\�D����D晸=t�)�9c?�~uf���������l�D���0��탻��wu!���.��!����s��mڸ��?}�:߽���N�(��`!wV�k�L2.>�"��}��M&�i�S��n�����ZjPZM��5�}����b�����6ot]��|���&�Ӈ�&! �p�a1v��ΓU4�|>룣c�<"�S�͕v����Am�z�DI�8�*h�f��v�p�;l�����3�]v`�b�8�v+��3Sn�9�.���&�Sô;���X��28��A�u"��K��Um�\ �so�ݫzzhE:l����$���P\16�D��3OOP�t�2�UJ��]K(n!�]Utx;���b��9�q�P�a�-i5n5�?��ׯ Nk��*�2���!�8UM�{f�R��ڣ�TV� @��""]]H�4%r��d)�$)
�������[�|�DR�qsF��B2�8E�u|>�^�V"�6sz.������ 	���$y� 
CV�	D%��ZLq+������<��mC�?	eK�� �%� pwF>��N&Yq�&&�8j);v��-Gyʊ��ݽ������/%څ.�9h̷B�ܿ~��L�EO8���������ٻ>]�Q�*H�p�ʉ��2�ػ�ד:�\E:l��]��ݦ"����o��]�$��1%�����&���;��뷧z��͞F����5&��nӈ��>g{�����j�^-�U��b���98��GH=3|$K���=���G��|'�A@Ant���;��ĵo�eթ<x�wo��K9�Y��O�M✮�goGĂh�I�fH�w:��,���0���ª1<�*������^˅6\�3MCL{���}��ϳ�l�X�p�t��ػ���|�\SD�D�md���mdc޻h��ՒΆ�*/۬ދ����D2�/��pó6�W]۷�j�54ݩ����'2uO�T�xE���P�0�R)�wV�-T"���N�F\ݾ�*�S�[w}��r{���Ba0X0�э�"Yy'���ݜw�8��9���U����M�m�`����0�J�����f���v��S&��P|���ɻ�%қ�DD��9����վ� ���*�SőTj��"��4�j���zE\�&�'��B�/�1%���B#P."�`��]��zK��W�or/%S;ݺ�ٞG.�uB32���]�S�F���J�v�w�RO=��Q��պ�����k�f��n��ݙ\<Ȼ-�zY����nG�Ҙ۲��t7�s�om���e,���v4d��Ey��e�flxN���tӻs�,��j^n�f�=�<��ݻ箢㇞�-��d0ܚ,�U�j9I�sG>݋������cz6���9R��9�-"vev�D�KL�n�nސ�k���ή���L혬M��m�ݷ�n�A4%)L�te��w�|��|���\�=C��p�<6R�&�����Vۍ���xo/�Wft�MM6�"�)�(%��<q�T����N������ٻg�gZ�ͅϐ+���Q8EJN)�g4Uw��7rwL��q����6�]��d��<�))��)\[�z��R�qyZ��w�}��r��M��Y3"�c�@ʆ$��@�x�>�W����v��wm�=����j��Lq��	�m"��7umb�QN�� [��ݳ�j�S�U�v����i��;u��00�F�K��Ӻٚ�EW\n}��b%�!.4:���	�¡�}�7���[�x�DR�qs���e�\�)�x���Kq�*M��ݶ�J�3y�AO.��%m7��z�(���UM)�6*X�/�Ge��`z8E��7�:b�
Ӝs��_2��i�����Ϸv���>���f�R",D��Dh�cb*=��E�|!7<���ێ�MM7r��_����ݵ����3L��8�!��[��x�y��H����G­]̾��-�pBJ��pn����}�֖�I˝];7f)������3*��R�I�LB	3�
i��M��T�|��W�hR�w�֖^I�rb]�$������)�5N�u��%�z�c9�^��>I����7!�h�$m$�S.1�=]Q��^i����j� 72sx]���e��D2�+�Q'tTW����>���n�K���ٻ8��s��M����eF����e]յ���M��sc���v-n����^(��1z��ut4�� �шsg�G������w���,��/_a�u����r����O�߇�g� B�zV��!�-�E=¯nZ�[�2v.*,h/I��qo�N�7��vi0��V��q�
L�~�{1�J���.�f�jq6i����2����Ԩ��:K΋\_>�6Q)�;���&=<�H��6��HQ�`z]�J�U=GU�ZH�9v����<w;����f!�Q,a�Fݪ��7b�@�Nb�O,��_�]�w���/i���x��gJ�eV)r�P=}������Jv���{�W��y�������+�Hr�B<��<�7R��8�����:��g�=��Z��� �b�|���Br
[���H+���+T�%�Ek�����
�����n1�uD���BX�̳���Nk,����D�\YO|w�t�tUx^'��^�\ޛ�m�3}hͦ�4xtӡ���3�<�{���mT��'Q˵�vΤ�]]����LmA�l�R6�^l>��Z�S|`៪رu�=i�ч�7��]�u��bI�R�i�qb&�D�����O	����FN`��.��s�Y���r$ьb<�1U�N{tʋ���+�(�����3�C�'wI�*���5y�ལ(��v��;�z��������Y'q��x#���v
��]�c&���"��o�xd0i�aհ�zBB�M��-�?[��xt[�n��[�)�J����D(�@��t"�,���=ǫv��A��*�A0/
���4{5� �0���B8�q4�����M�͂�8 ���˞�!1mMlW�e�R+��  �%�����;� �:sg2�3�0�a�����a�%̞��ֱ�:�^�n��ވ��&��=�H�X��D>�Ѥ�ӫH`vo�Đ�3a�N�@��K��k�)��tՠa0O�u "�a�^qƷ6q��ۧ"aR̒0�L�������HWs���#0t�<�W�ćV��\�a"i{Z���d����d� 0g����p��_�G���E�=��/��\Ͳh�>(��?�t˦R��U���<b�E�����֒��r��'��w��2����I觧��r�uh��G�O��,����T�
���2�#8����!Hp��%I��ph��
�\���s�g.]
�A%�����bE�F(������m%յh�t9.)������~� ��=;��<�
R��۸>��a�Q�>�:�a:��R)� � HF��kY�1h���9,����<z(��*c�wm��zw���X��,�{r�n?@�-�!�a�#,���p��PQ�q�'S��2���;!@����ݫr`K��.��u�5� ~[0�PD��B6��U&1�� �\!��F"\�K�a�oց�����l��?|�C
�d7���-�Q��7V ��r��j�Lcⳗ�m1i�Bң
"���i�Sl��cw����9/��J�*0�E���c&��܀M��L��3&'`L����4���i�W>.}�g�l�M��&h�a����q�cMa}@Q�+1�<�n�"�s��v���l���-1|�\���g���U������4$C��$�M�DLdb)�u�C�B��hY�|	��|��s���Z�1f��X>���n�hs�C^��
����$i"Yq�S���ɵ&�z�m��NE�b�,1��u6��T�J6��p���5]�|���g�3��:4�aU��s��x�I�$�s�-���5�L�ǻ�|�!!�6Rp]s�Y�f���iX�� ����Nj��76������d�1�XB�����}@
���_H:�Q��i��pj��Wh?��ˮ�����]Ѷgx�����s��}�����V0�!�}�u��I8�)��Ss�}�C0���׆����)1���n}���W+��ٶZm,�ן��<�ՊY
b�{}����ĝ����;$�v��l��w%xv"����Ժ�UI�Ed�j��m��d֚N�9��� �F����w�" �Q���	���&D(�h"(7�P������U}�j��ף�"RDbi�ᧈpՑ�핺���,خ��s�a��Z|�Nf��6�ͥ3��0����L�d���X��:��r/m�Y5�=��\�F���z;��x�M��< 	,$	�����Gu��_l��=�m��e��>��i�}������	>e}��i=�n���ٴ�^y��
���- �'#Jƚ�4�����ω&��`�;[�ѶV�m���u�n}����\�wf,�<@BO��`�{�x$�('#L�Ԏ	u�0�8����tm���ә��ox-<@d���1���J�aj��{�]p�5�!f���QN(���\Ljb|*����<���s���|���c�1f�i�]�����ϓL���!3���|���l�����t���f$��8���i}��Ս5��.��$����.q-��gk^6ɨi�!_>=w\�k�Y���Ll=~ͯ��V{4'�f'�;!�&�t^o�ԩ��OJ�4��������!�����d�w��\���܊��ˮ��_��K���Rx��;!;Y�s;6z��Q�mW\g��p\��7Sfc�[�(띏��w��;��8��>�u�O`��۳�r�mz��C�]�k
7 ����ޝ���t��2��p�V���+.6��^�]�E��q�Վz-��6j�#�s��+������\i��L�aУ�㷷[C�F��1���5�f��C�-�-n7j����:�g���@Gm�g?�v��ݷdD���]H R(4H �7wV�`�҅$"A��r�:3�C�7]��Ϸ������퇶��hu�W~w����筸�0�@�j@�tՑ�Wh?��×>M3�[;�7Fٝ��->�w�?S&	!9��&�����qf٤�.�s]��p�ÍF#)�a��k�B�}3���� ��|�&5ξ�Ͼ��|���c�1f�i��`�w�.q9$a$�9�k�ŧ��j�E���!����o�Ͼ�l�-�滼�m�} 2H|�k+}|��[>����k{�t�Ÿ��Q8L)F�{���U������pՑ�]��;���4Ͼ�l�l�fw�i�D���x�}�k�Y�xm�D�F	��q�cMaj�L���p�5�!g�Gq ߆��_`����u�n}��䶧�wB����5v��j�{��%�\C�<���L�n�B��1٪�P��6�bxfA�%�?=����~#iݍ �s��s�-����l��m���o�Ͼ�l�-�滼�x� |ͧ�ְr����f��,��6VC� ncMLB��g69Oن�;kq�[�T�x��v.v�Y��(��3]u���Eή���ݴY�w|?]��r,�}���ڋJ�bb��d��Ή2+,v�h�wѻ��T�c`�wv*!("�~Z�3	L�+ً6�M��}Ο\�4Ͼ�l�l�g�$���4�׺��ӑ*ciG�8���iw=��k�Wh��Ƿ>KOHNs)��֍��e9>�CHf�� ��EF����I�gYi�ĈIi����>�&ҙ�Ѫ4�X��}��.m)�N�0�l��揙�l�!}g��D�JG!Q�ن�H�ZD3��KF�I�S�����f�ɦ|��v��m��e&9Λ�'ɶ|��	����v�aF�F�t�v�'b��a(�eKӸ�{K.�-K�W������{�6�]
H�Mc��5�r����kH��w9�l�m��f���Č�&��[9�`�B0�!pw:��R6����6��r�ݖm�"CI�-1�����L�S=�5F���)>�\�.m:5@
��E�����*F���X�"�nͳI�Rs7��ͥ�iL�=�F�OzѠ�!�M����Lf{ռ@�S.�̨�����<�K�\F������7j���w6��E��p����F�k�S�ֹ��|ɮًy�ƨ�,�Af*#hKWڭ�j����oI>��5�C_v.豦��5��e��('#L��LK�#o���B�{�64��P������_�o3t��P������,֚]�(�e$�f��Ō5�P�9�S��ZD>� � �o�������|n��L�S;�24��P�UO������t�V�^qw:v�7M��
m6q�Yy�6��u���4~w��JY-�pBPM��q]p�k�CK��i6�O�|z��[6�ϳ�z �+MYj�S�u;�#�}}��a�(��Qf�i�Rc�黛|A$�k�Y��l80��ﳶ���kH��/�7cMz��GYg}��$$j1O4�sil�S9�h�L��)1[����Ӡ�6����x���I����m4ͥ�=Xz��&�!(��cM=��'��g(��J����b�?2��ݳy�����僴��J��2ț�-��y[�6�6#��_h��s��]���n��ogP4�'�b�<z�bʞ8�^�7Y���w��|����E X
M%s�lb79cQ�` xC��q�=��Tb��I�SK��N�����]���{�Re�`Ǐ��{���(�d�,��]95G� �y�eWe�m>�!����WmWi����×HHDfR
�q�_���d�gf%H5xW�? �>��ί�_�
t���`���`1�Q�&&^7��;�
�P��5v
T�_y*�V������²{���@ˆ��	8�T�z=U4����¨
埻��^7�@�[/�A�p�D�
b���|�+k��QԼ}�Y�&����B�U[���7i��H8�J(�l��4Ց����ۭ>:k�Y�@�@��f��M���weM�ٴ�c'|��������OOge��;����=˦�]��nv5������
;�"67#Ywc#�ͽc���r3�����#T��'Lf~��Z�*���\�p�n_u�=��D�A��f%��x�,��ۇ��������%��z+s��:���y*2<�.6�{mɭ�9��9��v�ŀ�У�n�9h��*cb�ez-��_5�X;�N8썻pnM�����|N��י�ј��y���[W/#�1)�g��>>�N�s��ƽ��u��O���ҽ������ #[���;/6:��Gv�6{5aE)"��H=t?��F�I�FJ�m��ΣX���4E�o��u����;le}�c7ks�utm�و�92�]2u?�ﵾ���3�hF����ww������*�Nq�Ss�|���--e&�I���w6�fҙ��q���#$��I�Zc����#i���^��%$F�v4�&�I�5֦�2I |ϒَk��l޷\��uZ��������i1gw�d�&Z���iC֑���k���M2����i: $�-��Y�i����:eikH����*F�����+U�ٶi6� �Zr���ϒٴ�s>�ѦRi�����76��`�ꪅ_�����Ϭ��"㉕��_6���l�fSL��D����Z�'��)����͛f�l��7׭ͥ�dC]��0�����c��D�箷Ht��W���� Q��IC�&DL@�� -Ij#H9`���c��5S�;�M3iL�{�i��e&7�;���I!�m�%���3F���)+���s3EP���f�H�ZD4�y�nZ��U�ۅ�1Z�/�{"�)�K�L���kZ���N�+u�G�OU9�݌L7.���a��{8`b�wd,i� ����j�xa$P�p�b�f��Up�sh-��PP��L���=����ٴ�{<�ѦRi�����76��@&��k���� ѐ&,i�#MD�=�w6��>Ke��f�3.�@6�O���>M�iL�/��l�4�e'���ۤ���#)�a��,��PT*���{kF�I�Rb�����i�Jg��h�L�0��*��;��^�"�=�<�'!(��cM24�#�gL�#Mi�
0��5�g6|�O�I�ߟ76�ͥ3��	�B0�#�U}�Kz���Ȅ��(�k�mۧ@�qp� ���j�]>��K-�;mg����UTv.�*1	R DE�c��k�C^ϱ��2�L����w6�fҙ�Ѫ<A$�e&�i�5֦�l�S;ҽ�J���AHSn7cMaj�}=7Z}@$��|��g�Z4�M2�����L�S=��Eg�D i6�O����g:F�f]ikH���24��R�l?������ː���@��չq�}1�-�g Fo�
��ѱ�}w��6�J��#&FOfY".*j���kg/���-��`	��Cn/H���Ή�pEmb���mwu�6�UckQQ�5X6��HL���w9���m��f�����m)���2cX�QXJ(�J�l������u�n|�fҙ��Yh�-4�Lo�wsi�m;  ��Y�6̦�I��JA6�֑���ir��v6�&�O�9Z����b��߆�5�P��?=����k������t��ʙnv�lzn����.غ�DO����r�y��7JeTdvFH�l��68j��Rc��M3iL�h�fSL����G� ��|��r���ͳI�R/��/(�`�$*2[0�ikH���F���i���ssi�m)�ϵ��2�L���ớNȲ$���,��:G�@���9	i��i�F��}�y���6��}|�sf٧�C�@!�i;���s�m)���h�)4�Lo�>9d�j6���H�[� * 
�z���m��e8��7si�m)�h֬�
�����L������B1���~Q�&6�6��L����?]L)��p].��\�]�u��V�{8(!��qY35��f,Cvl�:؉<�:w��(B��k�17�W�o9�m�o{��U�H&�0��*�j�h�#Z(�%����d,cE��6=T ��镄x֑)��T�G,8LQI�5�i�G���ikH�j�b���l��}ǹ���6��>�0a�#B=U_t��L��ҌF
`�6�1�׮�O]gk{s��n��Wg g���:��mA�
 +v��[���
F��1.�F�S=�5F���)1�����L�S1��س�#��|�Nf�����m)�~��La �p1L��5�P�9����(Ъ�5�,�<�Y1�}љx��v�<*�P5Y�o��N	A��76�fҙ�_}�6�&�I��q�����	'�l���(�)4�LW�{��L5�C\���7	��Q�j�����Zg���ϓL�S=�5F���)1�����L�t�I	l�5�bϙ��#��t@�����E'7Zhi�j�b���e� �&y���4Ϙ{栳Vh2>�|6�N��aM�w:/��J�Z��+^�� ⽛[��e�~�[�ݹ^�|���ԝ���(��ٝ۰��pHQoH$(=�*l((L�ߧXw�*+�Aۊw��S���y�l�ek���~�t��w�~�8�>1לu����v:/y@�����ȣƣ�T!FF]�55��e��"T��'�UeRKfu�R/J�>P½HQ|��G�~�ӗ}�ע4ems;y���a��/����n��N)���Z�6��Y�R�2i����YI��扺��:i���FK	./e�m"�y�F��[��������}A�W�"s��=3Ą�'b&�8n�dm�v��;Pn7�[�u�F�� �#���'��a=۬�r��B���5�u+f������C�����?v�p�k��n5�VƤ.����p�1Od���ӓx���N���w�f!Uӯ���x�{��K�t��^l�'�K��)~;��d�O;�BX�x��+2��7c.�q��r"k@��r4W,����xT_C�=V���y$`��ً�r���,������1�Er�׏�{�"4DF�@#s�݇��.j��Ġ�'iζ�r�]o���gI�w�ۏo�{���s3��m��=��������!�k^ۭu�B1%�謃Z���,ęcv=bs+4�Ӹ��9,��_,�8o���W��w�������o��c�g���.0i��
Y誚3��k����ET�J"�ʝ�K`�%��W}�k���pN��Q����\xctVK�Ļk{MP˾>Z������Oӽ���z|>�nz ����p����������Q8݆�����l�y�Vy:�O�����͵v�ҝ�T��s� ���l�w;�;\�'n���xs'#�v���v�u��[�N+�e��#�֞��=g�*�x��qt[�@�l���ce����������c�lX�]�n���3�����w��s��t�������"Ym�V���5��ݵ�t�l=�w%֜w���8à�7�ئ^8��8��]q�s��[�kq��=���q�t�:]���vn|��Ʀ�@���/
�Y�_X���:�pV҆�m�����b�F�F�%{]'M��	�K�m�y3ؙ�o��ks�a�{�kmy��=�Tp�b�5����x��>^7$�X���jl���Q�q��Noi�ĭ�3i���)Z�^��&�ٜx�7�`$L��[�=Tt��6;���L�����c��vx�\��7\�o����w;Z��;</Lܲs�we��Tn�h�ȏ�܁�*�w-�^HN ���Ŷ{c��X�FѮ9�6�l\L�ݜ��Zm�N붪�g;�U�ݮ�W-���;Q;��ɱ���n����Y̗omln���ө��Fϋ��+fL�9�m��v���!S��Y5��p��9��NM<;7��6���&���nu��Os��j��z�&���u����t��UۮƵ�1h&tq#�\&C��3ݍ�Hϧ�pu�gZ�c�yۺN�ju��'���P8��gg�k���u�I.W=��m���X�gf��A�筱�����T�s�yZظ��kls�s<��P<���/th�+��C��W��v���K���ݱ�{N�n�*�f�;A���u��lE�6�cnwݜ�u��8wkV�{	ۮar;/X�.6�\��,�7qU���ڼ0�79�켽
��W	��\�&,i�rv�٘�n�N];�Q�6��ly�n4�Z䇙��읹C�^��.<�]sPv���+��5��=���_�]ν�v9��r�Lc,n"�\p'Ξ�ė/ ���|י�xə��4��t��q�8�I��g�G#N5/������:���!h[�#�f6ޑ�}��_Q �-�!��DpQоE� k�^1�d���|��@�O#�g0�~�r"G��It�(�Am�*�4��E�!CH@����'�*F헏�t���}r��x�}��r�
 �](^dn N�g=� 0��:$�� ���^ߓ�g-�A��{x��	�X������r���� '�<�
:Z���!�4�择%w5��<1�6�T"J�^^�-`,0
�0ފ�e� `B��V����5;�Z�}�A7$��$7++i�%�L@$4w�f������*\an�V������I�0��(�2�f��ױ�;�%a�jX�mM�V������h�(RaXKnوD|a#v&!�8@?E��@kq�����|>�"[�z,Ʌ�V1���E�����3��ph�����7qkn݉��҇.6D9���ϦdI��M����6!U(�Ru#�P���D�+�6����椪[��0ݶN��d_5ݨF��H�f�Z���.�+\پ��9�{UVj��P�>��fR+�X`�M�kA��ʨ�e���4NDb���s[ѿRl��K��+,�À��b2�.�3�<� Fx��я�;�R�G%?K.��܁ 3L⒪�0���㝱|t?�\Li�}	,������:.�ޓ���ۦ�*�el������ـV�{nL�['^�q�z������ٱp��!�]ѽ��v���[m����5Hú��n�^�����FB˶]��佴b���8�q�3�6��nX��V���}VwH>�E�c:V��X��ۺ�m��i�-����Y�틘f�S�T�9;;O[OwW�qr[�r�	�v�ն;K%�~zݷ��lc[�T�nZ�Z1��V4Z5hٻ�s�5E%���D"ń��f�
QMK�a�H����㎝ �z0�v���v��S+���ԯU
�,1N0JQ8��H��dc��z6����Y�i�Su�q��� �A�C�C^��J�4�\��� �\�-\�i�a�Ws�-�����Rw�t���m2�z��a-�Lo|�ͧ@CMp��G��D�J�6����n��O��Ǜ�a��>�銆_2Hi����{s��6�����f�l2����S}Q%(�b]ik|*�( =��l����u���6��}|�sf٤�z�Ӛ���ϒٴ�w���ri�V�3T6m��e&+�=�ͦ��x�$'�Z�bͲ�e>�|n��m2�����L�5� w��MDarBD�Yc^W�:�]WR����x7�köXۮu?��{�Ȉ��P*��p�5�!����6m�M���c�ͥ�iL�7ѣĈBe����{��a��1��ό�TP�RREt!i���v�M���z_���V�fr.'��_Η�Zf�A����5&��.C毴j��S�*C9�t9��	q�~�����,�<��,b����q��5��C
���ld�2L1���$h��H�m5F5Dd�5$IQ�@QbLDa(�؂�h�4[���r�_�Q�cY~����i�G��s�jz@V@��G>�|������q��44�k�׆���e1�������l=��X�VG�B���ikH�����ۄ�9	i��i�F�P�*��!���u�i�Jf9}�sf٤�)+<�J�Kf��DKgծ�e&�I���cY���2Bڌ��֑���k�N�64Ց���#	 �;�|�g�L���fXe5�3�u����t� s�A%�^1ȣM�V�q\�v�����aLhn��l�(�gM�_��{����X���"������L���d���i)���h�)4�L}����A  |�g�l�kۦͲ�l���3�p��̒'.��5�C]��O�2!I�Zc��[�M3iL�/��l�4�e%g��M'�� CL�,�t��H9��cMB4�!w��u�a�"ߧv�C������Ѩ���FH�W��*�r�.�d��\ƞ�˯UJŃ�wp�osC�&g[�D��|��ҹԇ;����9uP�3_w[���V
,���UH!�zk���˒X�&�B6+&*���wjܢ�X�Ql�&"�h֊��Z�ͶځGw{���b�i��ϯ�[����V*�W6�}�da ������4̧��T�S4�x��C�	��BR}��Ҹha���A4ہ�bq�t)�[�2�Z�$�����2�)�s���L�W=��-4̧�'h�\g�Ṛ�k�'vq�l�.�+�`�q�J�p�f4�z�Ƙ�1f��w�{��t?}vw+�z���f��L�4�f�4i��e&>���m4ͥ3���,�� |�'̴�;��0֑x;�d�P��L���������� ���)�������L�}��m)�a�+�E��H��}�Gy
��(BR2]i��3_>�Ф�2��ܩ����bI&����fSL��9��S��>KgzzݩT�+4�ۊƚ�4�*����w��Y�Jg�~4�M2���M%�I]���w�7~��^Ok#�i��.t�l��=�B��V�L�s�^M�RS�	qO���qyR�ꝼ}���7*��i]��m��R�v�UEX�"�Y5�Qb�cI�IHm����H���jMh�ȰcF6�4�,�kZ,�-6�Nߕ�MUaj��c�\�[6����Q��I�[@�B<����4ϒ��_}�6�&�I�o���"��!�
��n	�MƓjL-�ƇCn3�Dƪ��yx67�����Cq��������]%�����2��Rc�uSIl�S7���Ͳ�l����!�H��ZF�`�0�#B�ī��
�����Mͦ���c�糛6�H��̴�5�b��L�S9��֫T����	�
����y�S(�"���Nj��)1�j���U�dֱ�M�Cv����;���䱯d\�z�%��P(�n+�#7�2��K�kýJM5���Z�����掃UT!��Yz���6�)��Ner�95�a6��/��&�e�Zeo���һ�I�z%Lް�|�q��9MQ��:����w7>�����d$��Vf�q�x��Y��,�q
��`�[���5`BEٌ]QG)JK{M�����L���g��������f^�.��ϧwC���������p���::�uq3���v�5��JK��%u��m����˩i^u�n#�x���Zɫp��R��cc��.�w�ܯuƇ)����y5��j�Tz�u�/�������l�&A�+r�r;���瓵��m�F�d��n6v�u��q�δ�+���"��-�b�۷+zz�������[�`�Dm�#�ɣF5EA�h�$Ƞ�	�/^���������.� ��n�5���(�����I�y|��Y.�!]�~�{�}}�&�):���->�B�(͙r�c������n�7g�SJ��A-��`��0�Mѥe���T3���n�|������`�^� ��]���@[�(d,�$e<�߽�ou�>Ю�*�g|�qc�N�wH�ZD59:�a*����1�����| ����s��l�-��}���=�Դ���$�)����a�e3�wn�d��*9$7A���s�<���6��@�{ة��f�}4�M2�;��U�CP
A�y��ci1�e��ns�R�Z�mE��S�f��E�>���o�{��y~��d�Vcg����2���1�j���e��xf�0�3�r���I@�3iL�;��ͳ	����,�،�E���f�5���}���Dl����=��D��D�I�q0(�g�y4S��.:gz��T�g��YQ��<��P�ѽ}\5.S�U�[�����xc�]t]�u�qϱ�)*�4H�F�F�VKE��}�ͫk��ޗz���ͦ�u�{�7�i�Rc��M'� ���5���:Ɇ#E(�Q��i�M����y���m)�_;�U�f_0|�KϽ��Kf���o�F�I�R.x}�"�9 �ʺ�,���
�l�w�|�M���i-�Jes�f�3)�쑐��r����L�S;�Ż�DA�3!I7/V�޹vk�!� 
��]6�M������i)����fڲ4�#� =��~8�PFXaR�)������QB�vդ�U˛����춋r����]���;$�2Bi'.�E�����80̦�I��\nm)�Jg��gUg����2ҳ�f��٤�s������a��5Cf�I�Rc�5SO@$�6�ϳ��Y�Zm���MT�[4���,�gd�Rm����^�VL�&G4�qT��S6��_}�U�fSl���*i.���<|�Q����:4�5\K�*}}3+����b܋(oh�tj4��̈������:2ͻjz�M�ؕ�J�터J�6l<���;h��="8 `�EE� TZ,o�E��q���˭�gɶRc�5T!�!�]��-��pX�VM� d��y�u6��%2��3F���)>����ҙ�쑁-����ϙ�ً�~�"X�EH��V�{8���TM2� 2y�u6�ͥ3���,�-6�L}�U4��%3�����+������<]���;sׯ�vϔUķ���m%p[�ϧ��T�-�)����YM�c�i��-;�ߛ�Jfҙ�_}�ٶi��-/=ǚ5$&�L�[>��h�)4�Lr���-!ME�ZE��!�?��; �|�Ls��i-�Jew�f�3)�R}�k�ͧ@g�l����\bI���F(����XF��)��+�i)���h�)�A�6�L}�u6��q��4Ց����}n��T�e���Kf�C�dL�{Fh�2�e'9Z�siL�?_=��sI��(z>����`���m��sg{6��8�{������Sok#�+��5����묉���}f"c�M��NT�YrVT�N�n���|���rn)Q�
D,�˻�0���;֞�5�CSg�����#�@c��f�I�Rc�:���j�C2W;�g̴����MT�[4�ʜ噣L�i��$������9@wH�&���qn�}�Y�sO	�N�>��U�\�+�nN�~{��_v_k�S9n|�g�L�/��l�4�e&+�Z�Kf����� $�-6�L}�U4��"���1��I�@��j��P����i�"I�m-�w�f�3)�Rs��Si�m)�����ͳ�&��Zs^�@Y����P�u�Y�"�߁�L��)7��&��I��}�{�ϙi�Rc�5]M����t�|�r��9��B8�4���@���w�W�Jf9}�sf٤�)1\z��[4� `�5ɝ5�!��!H�RCS��M3i_g��l��)���:n��ٴ�Q�ٚ4̦�I���Si�m*>�d�C���L�9�*��s[ܜŞˣv��;}s��th�p�����I�ia2�#R�ڃ�n�SQ���G�$�/y������r'�e�;=b��"��NN���5ہ-�P����;-�n{hCu��s��qup�=�lrp��\i۶�0=�����^�By��	/]\a�R:�va����m�r�V�kǐ�ob[���5���v��s���js�ܙt�ݱ�����q�Vc��ۇ
-uu�Y;����s���U�N8P!2���/KnS{Q��-p�qn���^{��=�n��u���	�~�d�
����!�m��۶��!f.��N���⌱�:�q�[\v������FvƄ)�V�~�PAԄA�!��ݎ��4�!N��4��%3y�e&�I[�s���I8�gL�}��6�M����}�D��l�ĺ�,֑A��pa� QI�Zc��[�M3iL�/��l�4�e&+�Z�OB f���{��ѕ��	a��5�P����Ӧ��k��걶[���2�麛Kf��G{fhѦF�/p���(�,@Z��if�KBd$0��]�sg��m����ji-�Jf�|4�M'd�!K�:��p֑/t����L�)��qX�VM��p�M%�IO�	;��l�m���5���L�S1���͛f�l��U~��%�Qh�YѴ�f$&S`[�JO[vMȁB��L�-���*��~{��s�7o���I$���\�k�5�P��:��i��s:�f䌁'��|�!}ђ��5�CJ}�})��P@Y	��i�F��/���/�r��{6�%�c�.C�F�F����'4���Au�'Z�G�?�8�U�zj�H��-�݅z��vfmi��ޣVA���1=�j�z+8������~�}u��k&��	2H�
��V�ޗ�ڿ��ٶi6�J�1Ʀ�٤�o7��Mx 
�F��9�y�F�QH[Q�Nnm4ͥ3���m��e&>᪚KO ��Y�ٚ6̦�I�s^nm4kH���YJI���Q(���XM��]ǚ�Kf���{��L��)+�q�M�ٴ�#	l�k�ş2�mB'Ӭ��1�$BC#(;�"�i�;�3F���)��<�~.|�g�L�/��l�4�e%g��SIl�S<�y�?�]��z-V��1]��ن��_n<.�}���������m���;�}�וֹK�7i�o�2������jm6ͥ3��;�6�M���?�i�m-�w�f�3)�Q�wn�F�1F��0֑\���zi�-9��<��i��s>�ѦRi�[����vH���%���`�s����n0X���5di�B�FJ�,�A��i����J�-nE9}=Ed���:X2�������=��Q �P1��&��l���jݽ��P|���3�q~y��;��x�.� #��؁L��cR�%Ǟ�W[�J�nN��`�(iUI{W0M��l�čۡu�v�E,>k��Va�em��w�&���8@:�)��;����F$�����
�8�b��z�w�ER�ݙxmT_�k�T{���=�=��uy�p�-�����������s\���遝�������vTl��u�*��A��٪(��/�u��NH���Q1WC�=�'&�;�՛��yg�3���j��]�L��(����D)�Q�κ�=A�r
�[�i#w�m[�w�}m�u=�E_J�L�Lտ�kE&�e<��"�C���*����~��{Q�i��f��yVT�O��{�����F��C;"У5��`u��ݾ��&-�;'�ŷ@^������x�g�������܊��/u�:����uZ���v�79I��ބIU�9��`^�e̅aȸ��+kL�Nn��IV������X$x�!8��U�H��v�:�VEL9�d�we�ָe9�������|2�h������<�;���#�n�:;��L>�X}�ޅy�w�g^IL�]�͕�f#z�N�$a]����\ҭx����wl��.�LR���ݔ�r���j�Z.��B���P3�2*�ōx6A	��F�*�H�u��;g�q�g�V-�	��|�{A�������#����N��V�\`�M9�r�e6�S���~��h��Q}�3U�=&�"m�y��o�����Ң�àh�9(2g#a;��L�;�؄��G�j�v�8p��-$�XU�8����A���T�­�:zy���$}��V1|�^�Waà��t+:�Nc�{���e��Jӕ�N���5n��,d~�ͨ��Hp�]�y<rn��n���;w�߉�
�S�H�(eNԺ�Sr	0�P.��#E��4V�-a*�M�.��4qY�D<��!R�M�^=9������4q-3�'�X��^dN�>ct� ��ӈ�D`"Vi|��\������z������0�Ǜ�ܐn���a�Q���2��~}v܃F-��������=�����n�2q�_�'�{s�A��ȹ��D�p%��h#��F���#�����A�9�9�uU�g�~BCԁ}�1�Ń7�n��&�$Y4BM���9�؍,�eP�d*$n�3s���@�I�n#�H�����(�t�N?�f���$�r�s�Z���{c�'��3l�>�o���9
�g�=��}��9��:,�z-�~(�l��ZN<�a� E'�
�B��M����0�׍3&8k/�0�j,�fQFN�t�/i�4��(��(�PA/p|����b�
���J�m��1I� ���4]r0�Oon�J�W�;�13&L��R�A;��9��@�кv3�r�+��'��i 
�g-����%y�v��}���w�~� V1�k�rȥF�HQ2?5{oK�~��6�fҙ����l�4�e'�ޚ�2�,($F"���"�o��Vk��&5I�RW�{����6�ϳ|�,�-6��T,��xr�a�"�b���qF�e(�B8�4��P����u�a�"P��<�}���4�2��O}��Kfҙ�{�`�P�dxU}Ϸ���l4
F�d�S�miӹ�	�׶�m���t\���=j�S~wi ��A$�.K��p�k�}�l��)1���ͦ���Q�ٚ=䘓�Z|�&9�카�6����n�RQ�	"��ݍ5�i�G.����U4ϒ���kF�I�RW�{����6���x�׀Ea5d{<A� -�e˛Kf�d���̰�sﹲ���2���2�r����M3)����0�=��%��4�3�l�)8��%�ϷW>L�iL�{�6m��e&;ޛ���.Z~��j�3ސ��g�W�iz����fN�������H���CĐ=�뉈TO�6�[���]ָ�q���1ѹ�������1�@hK�"$ETQOYӾњ4̦��.t�%5В, X��!��0֑c�糛�����9�}�%��ǭh�S�w��UͰ�e��W/�q�d|e�6Iۈ\���n��N۷<V��7�5�u%55D~kvn��Ƙ����{��ƙL{�*i-�a���-�a���排a��c��s��L�c��_5��Y��8�媸S4�x�Z-�-�?u�j�q2�g��Ͳ�l��{�w6�&��i_|�~��Z*3d$˱����1���ͦ�������l�4�H��ZsT�ع�[6��g�Z4�M2��sqΚa3��H�u�3[� T,�ݿpX�)6�Ls�7si�m�N�h�eB7�on�hi�y�����l)��8������i�nm-�g�s>�ѦS�~;���&Y������2�W칆ĕ�*\}��Dp]{�@���#��H����2*[N�*�6�[��2;�W=WPpb��8�sy{���*;�e�U�(�?ig{g.�d�
B�!�I2���\ރ����������>���[���G|��sm���m�^p�w�v�tpW`�tpu<lQ�y��;(�\���ӷP$tuljx1����4
�&kwh6�ڂ=��X������>�M�hi��[�C�w5�ΞLc�T�=g�I�7��'jHj�רJ�Ū7�=S�+��q�̋�"7gc&y�[�w>��rj�����m�d��D��h���_�L��^�9��;�����2�j�=9^{a�o6�8�16ێ������iz��V*�\�[6�'��4[2�)�}�76�i�c�~1�?�C�m��z�z��ٶ��>��ca��L�d��P�d>�54��iL���P�i�Lw�*i-�a�9�(�v �
J�9��cEVs����֚C4��]#z�;ճ�0��&�����Ri�����M%�IL����A&�q��qH,i�F�� j�=|�fҙ^�y�L��)1ϵ���L�v �����|�&�I�kƨJ)�`�F
l8���5�C\}�`�P�2�I�C7�����%3���he6�Ls�7a��6���w��b�F�2mlN�z@�dcN��x�F�gZԋ�����_��='�J*�H�+�w�z��B����i�3_;�ٴ4�e'�]�[� O�L�-f�4i��B���TNA"RA� i�>��p�lU�L�b��TF�
̚�XT�����٨�=?a��EVweB���qye������^f�׹J����f��*��p���X���UTAPT�_N�Y��}��M3iHW+�(�)4�8���fӲ�|����9M��E���NƐ3T#�^6�l�Rf�4iBФ�}ù�ZL����Y�2�O6��Q�M��&+.1��a�i��>%�^�M���=�����L�;���I��2`���q���Y�";�V�8Kġ,9���m
LW�;��M!���"s��ş!�����Ն�L2�w��L4�SĜ��y?�0�f�kd��Cr�Zv����^���Ӎ0k�ѡ��x�M�6�mlf��qT��ɖ{��f����)>��:�m-�JC�����i�-1_p�nm@�!�t��x H�(Si&౤M���M�m�)����ϱ�2�HRc��[�M!��W��h��>��-|3���KIF9ZE��!��j�B����0���}�;�<��xtp9$�I9�FDT�6�_fb�ukg���R蔸�8wlY��w�|�Q�#3R�c;-����o�lB���ME������-ބ�""��"�UUTETTI��e��E�A����6��0֑����	L�Uf��q�e�l��z@KL���s��Jf+��l�M���㭆�ٴ� E�=3����@�}���2ɍ)P� ��H��s�^���x
�u=���4ϒ��5�Q�Ri
Ls�q��N�@��ׂf2��"	�F(�RX����L�/M�M�]ûn�g��D@�pU=YXR�s��G�<�l"�i��}4�M!I���3g��h|��wעƚ{'_���b8��)���B�r�B�B0�߾������f=�����P�֯��%�G`�j���뛼�T*�� �������3+wv�%�0�EmBn���6{��=��]�\�32��dG�j�R��ک��j�]xe�T��\��%�{����)e�%A�u�@T"_j���'��T_:��f�^^9�R|�Y͂Xv	��q�[�6n�|�g�QV*����"i!)���mO�{���d�I�4�b����wv����O��Gs���c��^�}�D��F��5������jnCٴ>�r뷲��n�x�K��&�gc��=�ʚ�s�)o��q�)��UL�������ǀ�32c����d��5�[�H�-D��{�w���Q>��l�4�ٳhi6�N]{���p��T}� $��&��Sa��5�+76�CiL�}�����)1�t݆�I�>�K=^�e&���y��6� i��x�;R��$�F\v4��x%sd�f��a���tjKC)���6�Ci�D��V����=����B����4��vu�,�υ<����i�<��͚CL2����E@P��w�"+���ܜL3�6�j'��2H�
�WSYP�v!�JRT�1��ᱏu�s�˹0�],$?��:�A��Gz��I���1 $�8 �)+p1��v�N�܂���7����b�,q��n��ѷ���=vt�=p���j�\4>�[���PcNe.M���j�xCA��q�l�7��a=k���ݹ����8t76қ��&.6��݋<F���˱���-nl^�޷nQ�n�k%�TG�طF�Y�0n�M��g����Cq��ѫv�Iղ�ݶ�SM�D�	H$�i$�&�=�������ס��9鎒��sDc�G�]��`�a|�Ͳ�tqX�Gk��kg���v����C)���nm4��}��Hi�S�s��~$��>JC'}y�a-�>�z�s�����*�m4��<��͚O@h����r���Ϝ�*�s�ށZ��z	
E
l�ౄ4��`��P���j|�)1ϻ��ɤ4�ivϼ�i�P��=8�p�I+8�)��[7��-V�4m��B��Z�KCL7����!}�0N�>�8hi���O")��R7t&\����߈i����7�w����B)��(}�t2zri�TkF�\s�OF���V�N�m�\惚�Nb[g�t\��LiJ�������}���ct��[4�'��h��Y�����;u�aM���Z�F$-2�.8\R* ��(�OD�qM�#G�x�y�S}r��k?���x�ƖS��֧�Oa51x�xg�|��J��b���5�����JzhO��U��}���t�B��0�5%ș@(& ̒�5�E���jKC)�{榒�����f�=UX�B';�_�nD؎ ��F%�����vy��>=��{B���]�/;!��)9u�y��[6��g�3ܮj��R@P-�����G� �!��*V������f��M����������(2,���{}%�0H�h��������w6i0������a��(w5ѣ�Ri
LW�q�ͦ��Q�Я�临�q�I@ى�؅�+yӶ�N�6�ݜ�-��/a�^`-k��1ec���`�� Y5�� �4֑HQ��h�)4�'3��g�ɤ>`�yy���}�#�m�Ә��l6�C��OJM!I�s�M���c���!l2����4����;Pc]e���ф����4������p|vx�pD��"�Q9�I�������_J��w1��C6w&�Vk��݈J5�J�d��U�Vо3B���~�d��G��gI �I�$̂P�bF�f��I1)�_�ܾ��~w��ikH�;�3&:�.s�Q9��G4f��Ho��+������I����l�Rr��4�M3Ѓi�^�����C_wċڐ���@�R9� bm��f����[6���'�]�SHe7�����a�9~l��)�w��1���e�#�����M\��a;u�;ix[�t�2-۶\/bxd��t�8���mvm�e\����ɔ2v��8�M!Iϫ\nm)�3�w9��`6�2ә��lE��!��:�l�h�0�Ɵ����+��ᙓ���w6��.�����L�����Q.�p"��ZD4�~�sf٤�Wپ=tKO@���uѣl������M���S=�X���8��\g.1Tٴ-6�-9�P|�3iHQ��h�)4�'>�q���6��l���_�bӇL����)�Վ�x���E�Y�T���W͋P��k��ʪʧ4!J�Qk�nLse	Z+t�ő�����=�#���{�w�������� ��%@D �I����`"f�?7�s�7c�4�zz�r)H�[0�m��(}���2��_H<�zT�>`s��6i����.�Za9�w�.*8���v oO\Y�Tj&Dn.:ݶ���m̺L��0�{۝��{��Bӹ�}sihm���s�4��e>���������k�P�ZM��E�� djT*&.�� i������< a���+1��ӮPdY�}�i�X��W��RHĄ���'#v0�0��/��6�i��5����HRs���4���˷�ch27���Jr�j1-��47�T�	�~R�"�Ng��������b�B�������8hi���̗"M9 l�`�2�C)�w�M���='��;^ޛ6���}Κ��k8��1P�n\�︊� �SnW��:k�։q�N�0��b��WrM8�W��7~=vɑ�k����|�F��)���i���;o���ӧp��m,�q���-����8��I�8�Ł��5�ɥ�N�{f#�w|�՛Xӽ�LQ�k~s��6w����i�R�Y��0��a��$Q���e�Tu!=m!�7��l뼁kN����D�|D:��K.���n�K��:�e���¦m����FIDh�rd��9��X���O:��'��A�1�mfʛ��릯zojԱ�Kj�U�953�a���S�z>ry�fG�T�}��y��T�~�_J�ov����k��J%=��8|78�4��0��ܝDu��i�3aRM�/ox��>��p�=���Gg�򣯉�����7nz6�'q}�mE�����jї�$7��Pw�UF���Z��	Cvn�el����B�M0�nN��1Jd��t�P����n贿 D~˱��Ih�nD>>���oj���\㾣��M�b�4��7�ޱ�q��~�/��A�ڏ�p��F�u�p�n{�]Ah�꺳�1���8GC��ه��]K}��,1D�pSMw���W�8�'.=�0� �Z��f�!OVd�+WoE��������?OH��pb�8�]���P���=7�i����Z��a��RvWҸEiW�����ce?�q�����uD���
�!sQدqb�֭D�s�Cƶ�닺�ʊ���Ӂ�f&0o{9I�n����"GwY�ȇI���n ������"iI��i� �y�qk.��K��9�@(	�Xm(��A$�r�q{rݚi����q�:-����Ws�n��ضٌC`�+���c^�t�ۍ��p��t�fr���{8���۟;��:5ؑ����Et<�H�'������6{mE�k\%ö���#�Ymb����km�9s�qգ�;{����S��S��t�[k��kֶ����m&:Nz�cL�[Pi��æ�W��!��y�S��:�uDv�n����n;pcd�g��uܛ��^ٲ��%��=s�Ե��ӓrc!�Y�=>����7�e�Ps[�9��N-��=)ɸݥ��>X`�%.�ћ���m�[���;���<�ǂ�%�']���Y0[�ۛqU�ғ�ڗ����8��.)4u!���u�j�5�����u����S��M�:��9�
��J�t��7V7N�y�d���\��<�.��}<vUc�ޘ:���#:�9����B�8�A%��
�\Xt�x;\p{3[�eM�=rN���\9K�zի��ם�d�y�9�j�걙=�;�f���99.ɕ�z�퀙f���ۓ�Z�]�;/���N�e����Rמu;K��q��oc<�cqs��^�<�݋�\[���]]F���Q�] ��w;��*$�����݈���ȴR���4d��&�{pnƎo��*m�ݮg��Ȧ�V�RWXv�w']Qs���ŷ=:�vw\�]���SۉήV��v�\ڹݻ;\�ы��U��3��u�vmY{^ |w=u��k�-���a��ǅi̜�����������ۋ�"���^`ƞް\�dۧ�&/,���;f���n�+��O�{Q����Bz6un���&��m���Qݲ�w>.��s�88�\sv���#u����.���T�����'�O`��M�un�n^-姆0�F��ݙ5;ԅA��m㳸.�MN��Vu�m�����{^{39����^ۮh���]�{��`^Wz��_j�88�j��2�Rp]>$ӎ0����li=�T�:���\��v6�����`��##�ӱzkN��WY0�{�&o
-T���`�z�{q �.�A�0T�HR�;��C1��@B�S@�
��C��nqe�=�Ăܣpv�0b���� ���#�d�#��q͑iv�g�� �����3��*�S�g����wv�=4xN,f���w��p�wE[�dONaY��{|���+I�c��P!�e5�Z�<P�n?x�f�͢s���ǀ[ᥳ��#h�sb���J���Y�*D���ޓ��%����Y��Mܣ�Z�q��@X��,���=4@˞��e�u����#�F��Wf&9���`c����!7�;�10�H�{��om�1�-��6�QY)'V=)Š��rBJ���ڂa�DDwT���"�R��L=&!��1s�̓_^]M�$���gt�E B��o�'�8��us��j��Jմ�&f\����a���iV�]��= ���/����� Ǟ�@O��)#p�-ӓ%��]ELq���.]�DI���Tt{����������iw��'��y��9Ё����u�W�*A��ت33@Û:������)�9�ځ������g���wf��s�ҿj���׽�����&�������6���Z�i�tޑ�;�S��t���1��<hm����ϩ�la9���7������+Ɖ�p���GI�Y^�\�V7e���Ip\d����H�.��s=3��t��v�6�ɺ݄���-�ۍn�;�Mˈ��N
�gcv%]u�{e��K�OWg���)�(rl�n݇F��uS�LPk��g�<#v��@�ڊ�ϫ�u�w�yz�_,S%d�M>��I��2)�wrQ�N�߿�_<��^y��-K�����9��&���sF���v��6v@�w\�c24[��F	M(���V�d'���ݰ�kw���l�q�{kG�������V��4��ۈ&�n0P��Sf��N�Λ���!�R��J�R��s?w�6���<�cZ�5�Q�F��j2Ҁ�m�a�4����֡��2�}��M���s�����}���lv����r3��
�\2�O@�=�s��`���Qh[��<l6�i��/!�����Y����D܊5 u��H���{E�CL2�@ǹ���&P�k�*KC)���\�i��!^���LP�u� ���l���X�1b�[���'��]ѣ�=t]���V�8�j�g�l�E0~vжO�}|�m��(}���2��S��G���%3�Y�4�)�����`��(�ZLKM!�ӬJ}}mc�٣��lU��lӜ��e?�+ڡv���U��=��켾��؊
��3��n�`#N���`�SS�� v�u�E��f�b��}�Z�EDDF$DE!���%�2#bUQ��/L!�ƾ��m4���b��Q�-�S_;��i�>JC��:l�h�0�&�20���{㫛L!���4��Bq��^0{����|�C=�d�e-�5��8a[!�JK�#��)�(0����w��m2����C)l� �g��[�#i�}�m�H�QG��ౄ42��MPi��)�����e6�S�si�6��{E�l�$;�`陼�m���Z�1��v�:v�l��8��E���=n�a�\��N-�S+[�;e����7��>�jKC	�������:�����6�(5^��,�"�A>�S��cY.M!�Ǿ�l= t��=���-�﫝�a�L!�z֡�i��ސYF�Bܐ�|F4�?w�,a��v�E� `�#pّ:O�n^WgY��:|9��6I��#���(�`�x�N��+D�wb�wUl�5��*,>�_������^|,����> �`_M�e,Rbf"�ibgwD�(�i#��N����%He1�������撑�E���5cYڀ����0�egִ�S}���H�ZGj���}�m{�Y^%8#n4���S�H�P�ȳL����}ۮ�|��}�4�0�}�uԹ�L��{������Ӛz���.yu�3��l��#p;Y�n��6{qݟ^�t�q��=�j��Y�eu�ٔ�{�76�f�?s�,�4�)���ݞ ~a�S9U���)�uX�p����rE%֑���/�y��zH�aI�{~K��egֵ��d.s��#���8h_��ۈ&�n0P��,aW��]P$o:��
�I����i��y�f�00��K{����H�ےtx d�A����g�Q���* ��*�<d�,���m��\,�i>��:QtE��c�gZ��L��rv�glIf��;��)����3"�W^lp�36y�ơ��7�"E}����+��L	��1���$L4;�]� ���i2EE�cX��2��`�@DldߜB�b큦���}ږY^e�"n�-8��da���wo��P)�|�N}���f4�@]��q?U��ڑe�c;��2�WOgi�7=n9&,ci+�޺�f�}��p�m9I�"j7F('/����3�e;�w���P���(�FRiB�>�֑�4>��3*B��D�qD��4���}�5԰��@�q-wK�e)�9����a�=�iBiP�s�<|DS��i�`i��2U{C)he1��˛M3�G�s��D4���, k\���E���\HQ��i=!�-+���M!�}~l�a��y�n�i<@���b���Q߉�X�0�1Iˬ#��(,�a�#����L!�u�2��{�����;W�Y�5Eŗ��v7F��.߮uoq�vo,O�7B�Qxj�ܯ`��
Fm�q9O�A���m�����at�;�/�.����Ym��0�I�knM[�㊍����&:����^�����Q�q��;��oS�=]iht/^�I����d����l�8:�8�hyh�n�ح���6�A�7kn�3=z���w;z0��v�q<Y�նnݦsuE�՛�{i�q�gܝr#���N�c����<����t�9Сò>xn=���6��oZ���X��r����~��(�H��PTE�I��� �E�ؒ��(�lI"� Q"��R�b�2DK.�ą#y�v<�hu��f-lR�u�Nն:��m�r	�H(��(�R4#}ޜ�Ho��T2��x�ܳ�3i�>`��l�G�x�?2�nB�@� �4��Ĥ1�\�$�Ф�����m��_�4��e;��݆�Č�)r��
HJm�$��f�20�����]iCl��Qh[� �R}�;A�0z�b�
n� ��m�M��YʪT;~l�O2����m4ͥ!���V������u�!H�����FG1��Պ�a�G�큤Y� x
!N�%��aI_}Ǖs�L����Zi�#�
~���M���ST�hD�Q.Ӷ�j�q�ܝ�c����Wg8E�]�[�W4��n�$Y�H��8E��@�������Hf�~�(��M2�y�{a��m)
�:g�Bl�SL�Kd��q���E;��U����S�z�;���p��hM\-�1��F.���N���5ndf7}
��ۘC���UIO�3:vwkt[W����鼿lŻ�޹�k9*(�,����c��EE��-d�iE��QQ��,�
�Y6+(=hw-�[w��m+���i�JC�'Tk�@Z@�/��0�M(ᚪ.m)�3�b�!i�Ro7�0X4�#���O�agAce�7���d�|���m�`����
�W��y&H|v���_X�y��<�񻥚&�$K1�($�"�.�D�}�wz6ow��T���Wiz������		iʉ���Ѻ�p'n#�ۮ�۟^{n�QGA�M^o2jm��f"��^�J�<�UJ�i�m����w��Sa�_C-©����|>n3�.��0�ʕ�ݱ| �}�6R�
e��:Y��wv��]�=�G�kVNC.�κ��Q�v5�$�-G*���K4�1@-pZ����-��׽�..��}k*sG�{���:���w�8�G$�';�X	�ƭ��Ek@clh�Xض5zV�*ش$�}{�/wY����͟w!��$�.L�n�� ;B}f��u
T�Ӥ�g��B����߻��h(�1�Bn�n�*�^ o_�2���U)[�������ڈ���1#��z�u�[�X7�X�l"l!��^\���I��>�^x�A���7j=�j��6�I7�;��9�	���%� ��$��n.�B�|�i��J�ں�*Y��j�ށ���^���PI0��D�M%����w�.�h�����fZ��\�ksH-�a%��L+W|>���bխ��5T�6�U�<5���Pg	�{�&K�ܸ�8�G^H�}j��5��;ۖ�܈��pͧ�x"2�Nj�����ٚ=w�;��2�{td�ͭ�����أPZ5�mQ��h֊����j�M�V0R��FKfR�}��Y��8Ȋ&d���}Ͻ�ƑZi�UQs�1D�i2��]Ƴf�{��E�%$�:Fhs��(A)Q.C#I�$0�LN [W'��)t�m��0$�..u��v�Us5��f�XjFcKF�\4����a�!�5�1l�ZL�7Vz@v����w�,�M�$/�ex�m�B#j@�U��}��>�JM��3ݗ4��,���b�"��#y�+�P�ZD u����r(ӎ&��!cM24�}�ˬ!�L����7<+�����]���j4��)�Ϯ&�E���Au�Y���k�Υ��2�s�(�f�(c�3)L�)�n����>}��ۉ�ԑ�N8Y��fSW:b�l�e<>���f�i;�wE�%��7��1F�i�Os�����\z#�,?uƋ��y�=��]F��ߌ�����y��!t�wn�55�)�pB��B�Ttn�uu]Dn4�YӴ�ʘ\x�f2��2�pb "YB�4�p�n^�	�mOd�v�p�a�ȼ1Ї<8�:ˎJ0��7&�v�zB\l챀�n��\v;tCE�fK�A8e�6�{6����2t�eW,�=i5�V�6$�n�t#�q�.c����ɴ���9���mJ����A�P��A�vԶ�ǹ7[�=7���F��z.�n��Ե�F�ۖũ���Ź����<Ć^�nq��*�Z*ư���,��/ҮF�EE-���E�MQ����ߟo�sNcY,�ୗ�	�c�8^��R�wVz�u�sk��k�Ynt���"��c¬����4ȄS��r�)2Ͼ�Y�8�s$����Ha���}旓JI�GiE,i��Oc����0ɋf~�;��\�=p�8`�^� �3y|�9RD��T	�s��4�&>��,��$v��wػ6� {��� k�t��H�0��.9��L��福f�=0e�@Ưn�� wU���x,���l�S�Cq���E�٤��;��L�'���l��3��}��fs�M3I=w����E�N�k�I����v񹘚�^x�n˰�9ׂ���*2p]h���ߝ�o;����|�\�e&Y߹ݖm&ٔ��Θ��4���6���ﱫ6�iuF���!Jbӂ�B)߹�]� �Woy�Ă�s�ةh)�Wٵ>Պ�>��sy*�ˬy�p�]��*�v�R&�7UsA��:,�ۊ/`uS�Q��F�}D�1cI��"-��d�Fъ�؂�#"��q�[!͸)�$Y�n]��3^�[^q0��$�i:�i6��{�Ka�7�w�~$>�w�.���w����+M�{j&pB�U��l��L��uɦ�}���L3��f�m= bg���Hi�]��!?�l�D˱���G����dVB'��}�>I�s��D�C_q�lhz����L�L�ܑ�b*�U��qY����yܙ!�@4����6ra{:���4"��2�4�s���44�<t+��a��^Q��6��;e�,����rH�"�R8��˲��Q�@o�rS ��<��Y��x �`��q�N�P&�1F�*����j�>��\-���q"�z�����n{<�w]Z����j:?=��!W�6�w ���{+���Q>${�n!���J�
���gul�xnݗO�0+\/d��wv��d��7V�Uy[�[u���~Ƈ4z27Vy�έ����i\i�nuӯ����4�V�.C���s��q�Fit��E}
n��vZ:d��^�u��zw��M�>��ix}�<]<�X���~Ө�nv_l��<��v����h�<��[_�~x8w���<ٌv�&J�8�Gj"T��-�c:�D�Ǽ��LB|�Б���f	��6�TS�&C}�棻[욿��$w��>��Ǉ�,I�|q���� ��ۍ����>#�.�����d��o�[���!�\\ʄ�v#[�7�4��mp��{C��g�ds�b�1��T���4�ҦwO����bQ�����r��Ί�ΛPun�:gl�����Sю�ȷ�rh还����{����tM~U� ,}/g�{�����}���.��V��9(���g,��b�%:�6�F����uzJp%�G+}L���=�ck�>�G,T�ܫV��9�u��3h�Q
d�݃g6l�F�h$���'%4u�k�K*�hh��y{.-mF,6�V��b=&�f��?o�뷹��U��ѦoeVs��ز�$Ǝ'�f�5����t�F��=��vOrՊ���Nv�	��J*�S����m���Ĩ��ʗN�ky���h;�� Yt�=����5�)�,l�أ? ��f�wNZ�On[	8��<���ԏ��OZ�ܒBҋ��]ù�i���d����cPTخ��[��K�}�1�p1��{��F�h˲�N]�����7�������50�.((<z��g-�'͘N#�"�3JI���ۣ�G偧�G��$
u��J�(ye�. ���$���1[�����"[C(Mp�i����H�P^���t��n*������ku�f�`�+vr*6+QDl�ҕVB��3B�GW�C��*#0f�E�ˍ�q��a��Q�e5"s
J��8��q熷�];�|2�L�c$�m��6�P�*,#�l���B�=սq�^ߥ�/x���;y�gL�Q��:�
BoW�W���z\Z��ٹ����ٴ��[��]�&�N��v�.(�S:~k&��FV+�{J�4��o��Cpi��l�9(���bx�����Z��P����˫\ÚzȰ*o�<p�����xw�Ps[�{^���]�,���5�&�$��T�:Z�i�(�rJ��Ŕ��Y�/��+��g��<��܇�!U)]U�'+]�4�@(���Me}�1����簎���`+H{ޒ�C���)v���#�4�y����]ؠ��<�m��v�&��z�7��=�Foq"�*�e�������Ս]#r�"�o2�Q����V)R�^��9��M��Wr��.wy}}����$��r�}��dD�($��Ë�m��Q�H�x�W,�E~�gz5��8�4�yhW��2}�9F��_9��U`� �KclQF�*6mL�2)H�a����6�l}��i�;ߺg�K�6�q4S��cM#�(����T{���&�?}ΖKa���h� ��v�����H.�[��� �8�;�Ka�7ι-�����up�)�
����y0�m�a�2&�I�s�P��mS�kE�۰�"m���^�f���!1#P��`����]P$�O҉o�Y�D'��}��������<��YɌf�7$��s<B!i9��n�I�{���4��@���X�
�T{_y��҆H�D�X�CH����в)���a����d�C|��ZGW�' �H�B���"�(�{�﯄`�>�a�;ל�L4��z�<�{z�o��S�յX�nv㭄�˖�:T�r�LG�>�'2��0ЋZ�L�Q]���Ι�&��[�_�>� D F�5QE1Y��4�2F1�����~�t,�F��zI��D�H�q��x8��s��d�O &��&�i&>����	0�o���I��{�n_�i�b�S�õ�pHJ�^�[��f��]���<Y�]-��\���v��9Еc���=����a��ݮ�I�s��sg�>B�h���.�����	AD��������[���wc��d�������~�&�)�0Q��)�����3߾b��|*d��}~؄���-�IJ���g�VZ^������*�@>���̽��!��p�k�Bd��3��0m8���z�Ʈ�3$���0�*|�;��2竲Ŝ�mК�̍����'r�NU������隗���ë�n�Rq6�����c*z^�q֬��9A5��}Ҵ��4J��0� ��:���Г�<�rq��ǔǮ3`�us��v�N��6��;Ѷ�gm����s�.��؜�o96���#��+n�n{WI�Lr�'!�u��v}�nI��޲\�&$�^:���v��'f�rs̾:�ދ�c�;�'��^��8籰`�7j�j�92]��%����k��ns�]��ݘ��F$���A�$q9��$ �4	ѦI�K���4L	n���y�;�x�9����c	��s�F��B�|&�j��M����\�Ѐ�
$�N�m%*�R_���x�;�ܮ�b�"|�{ª��H���h�Y	�������ޟ�����W��=��Q���A�T&���L��x��wp�}����7;ު���IP8cn+�
{�^��=��g���Y�����{|�Cm�l�6Ȫ����<>�3}������]U���#�n$��鱜6�Su��s8�U�d�d3϶���Z�e��S�'!a�L@�R#$7����j�o�fc�x ����=�� �h��m�M:���f��k5{�)��V~f�UJ;4vv�M�({�����\@SQ!����)
/
��<��F�������;5Q83iʫ�4��v7�"" D|dd`D��@L,�Ub+�����w������UV�í0�+�DK�܋,��	��s��g{�C��31z29#��l��4�y����z�p���`�w��©o���߻;���(I,����z�p���jc=����1� ��/���!��Ԁ�IӺ�#��-p��:�q��p�]w7 ���t�E#1�I��b*��*C�9���⳸L�fƿ���W{�xB.!?�I��6fb�;�x /;�蘽��U��>.w��AFa��0����p�sw�O��c��f��/-���f=����::��ɬ�y�W^J����N��6Q�q1ؓݺr��=aE�r�t(���|��_W�^�h��,b�F����hѢ�������{�3����(�<�Q�e �w��g��=F����|�n�*����ܥ �"�ne�߽ՙ��+������޿n��{㻚��{��(�d2z�=��yNp�7�jq��=�v�eu�g��F�t!!��)2E�����>7b���]��3����)A,0R)�1Y��|*�n�L߽�3����	5{��-!��e�C;ޙ�݉�}��w!�s�GU-9��m��)�ӊ����}��<�!�n�Ͼ�yFW��c:�B)ʖ=y�
{�O펭q]|!��:ܤ���d?�D��1��Jc}�g�{�FY�ҍ>���M�I��t7��5Tc痪q��yёQb�T
"-2#EF��66��_=�j�A�0�E��P�hUIŝ�UUW��x��{�������-h�>������UT��6���j���r���1��u���rv�)��H�bIn����ݣ�}�4/4O��U,Y܅Q=���8�Pa�-�Q��� ^G��u$��l������oŵa$�@�R�#7�̓Y�N����]F7��SW��PB��2!i$�5S��x�wzɊ�mMp3xUI��*i��M��m
����>���z.o<}�U&��3$j5Q"5��ALU�7�ɚ���3&��|�}�t�[Oy]��ڹ{_!���m�_KYիU�]��չb��nN��يp���Q4����u�e7	A �,�a�a��n�v5[�j�of6-cn��9�*�pOf�֞,�{8�s�8㛛^�t���t"rM���Cll���=���i��F:�WgJv�Ĭkz�*�vNv};BׯcpI�plݹb^�p{'/N�`I��8�ƚlg��c�y�({�U��ˌt{Os����î#\��ҋ�=���<:u����y�u��c=��� �t/K��m���j
�Ɋ,AE@�"(B���"2�d)Ex,�%>W@ko]�[n�,H���W/�uܻuX��m�m��e}��c��T/��b�;����}��㘾�I>�-���q'M_�U�>����'w�L���� ^���-B\��h��pnb���㘾��Ӟ�Z�{���|�-s��Z	AD�Q��؊� ]ޅRb�z���xUW��c�E���`��!�KF7w���{ϫ۶���n���]���z�E��L��a�`�^�`l�y�Nx6ݻ<��r�Y��Z����� M���$KeI����eYǢ��l� R���S^�^�D�p[be�M��zg��=�6�]��_�~5�)qT��w����]��A�#�J��r=��k$��Y8�A����.�k�oK�]c����n�����&4Q�4flQcA��d,[]߯_o=__nEnh�}^ݞ���(�,0R)�T{�"d�^i�������rs�l�f
�M2���!�T*�|�o�sC=�Tmgr^ ��a�����l4�e2��|�_|>��3���D��|0g8\H�bz!99���T j�#���vP���vY�R�	\]��ᄢ�������=���=�1uxwﾺ����T���G�i��)�C�'pr��
���47���ů������� � ��(�$)����SW�U7�\�����Q�ѯ���.�)9��U��Yy�����̧TaA���}������z��3���Xf��ϰ�j.�}�`�lco�u��h�M�m�Ɗ�VFԚ�D�	���.�/�9٘����m�#q�I�S^��s��*��c'�|��*�燚PB���i$ӧF4"��stq�}���k?{�y���x�x ]&9Ӈn�6�\��wF�ۜ�\z�ϭN^.SEW���[2��8Ñ��&�ޱw���*�������}��<�j�Ek��	6�
I��Fw�W��U��w�]Zֽ�)����Uc��gL"6"��(�y����LG�UD��7G����nl�_��h@��@�d���������Ff(Y�UM_����vlE�v�l5 ԋ7v �vM:'�mT詸�*j�[�nyd�����v�[ԧ��u43����L��l�V>�m�Ӈw��l��6�f��ֽ65���m�j,k4�+fX��F��DH�+����~�o���QM`��&)ҥotr���>;޻��	�����1��x_z�26h�`R'!��{h�R�œ�c�v�&_���g��Y��r͸[ru���D8DLn��~�SJ�o]ͬ=���&Ͼ{�ϻ`�@��IH�lS��*�>���)���
�P�6u 3gz'�@�$�I-�m��z��ǘ5]�c�ޱn�o�*��[� �%%�
E���^��P�zQ����mOo{�H���I"17 �w^�
t� }빵�q�K6}T��5:f3sν��\IA@�g�vZ�ˊ��)SzmN�(�u����l�bl�򷓜Ԫ�d�	����c����RC��Ul�ɼ�j�9u�*Vu��s3^�Yf� �Eۻ��Ż�y��d���}��,g�^`Z�{�4���)Q��X����wl
�Ų�p�N�F�XCĶxo������|ǔ.�^�_���X�`�?'���{r��4�4�C9�q��	�(u�Нz�̩֢�7:V��ss/XoE&��U�+ DƬ7b)!5jr�9VU|_;]�Q2��;�[W�Ag�
C%m8�U���,�2ų��S_MW�����6�\������+vW��[�P�T�߯%N����0���˫fB���ɗ9H�\h���֜"-�q�q���Ò�����Vn��3q�1f�����"���6\;P�3��0k����8U���p����e6�W=���6ޛ�	JX�?{����dQG�
6�D�=�6�T����8Y�����K���{B���#ˏk}n��o,+;0�)�<�tM�-Ѭ�7���L�۝�{�\���)ޘJ��]$��f^�K����zPOp��;�NEb�rw:{v(dr�@�ؚh���;��Wg,8%�t��b��K�d,�ѭ;�vڜ�iѱ�
�ӒD���]��B�B�� �3�[���!����&��5K��B��x��v��f���c�O�u�0���7�W�4�
�j&�*���<ށ�ovzc��V���}�`�7���/U2#�.z���q�8���q��b�����sxosy���]�x����G�{w�ɫ�'��'Mă�������Of��z��m��ێ�e� kLm�[���q���g�/"ez"ܖ�{G$�.2ݟm�k������3g�}H�ۍ��˝xz1�]������3�s��W�n��\�z���M��3Ƶ�v���=��"x��hKv�l��n�t�SS�ٕ��h�Y��[s͖
�piϕ�\��+ڞ��u�\tanN�^��{<nX�rn2Ŭ�x.
2��69�ݞ��\K�����u[�\<�3%���E�8���v�/ck��8&˵'+�獍�=l�
e����nyS���:��� <�\1���;E��Wgku��A��av�sm�Fk�K6��';Z.3s�)n�1���\�+��p]zx����nzw�c���{;u���v����'@�g�8���N�8m�s��`4urqOt�c���WF)mќ0��A���[��F���t�r�s�6�!�.����0�(��c;��M�����E�x]��\�s�a��n���q]�d�onp��u�ˇ��4���Zݮs��w=&�M��8Mu�`�6�״h�[q�u��׀�`��A�.ɥ��d�E�n�����ػV\ک,q�p��-s����m�hsrm�x֞��fݵ���,�r
t�q��n;�\�;a�u�.YI��Ϻ�l��r�\݂ی�l�z:x<���J<��s��q����y'�V�8��n�kt���%
�e��d���+��i��(�;z���6\<������R!�P���t8����Z6���xOC���\�7����ϗ�Y��l�������&�6���U^=��V�d��J���x�ϱh��:�6����&��e�0m�o,�t�<�9-�Q�nϖ�"wY��]c��;HC��4���YGCm���×F�l�Ml�[f�Kn:�5s�:�/oN��	sW�4<�/hŞz�ź��;\�9ݹ�z$��fn�񃮉@�H&�����]�tŠ�N��0����'�.��.�Qx�pr�qs� 7��Et��݆�m:L#S�ׇ7�F�;�i_p�פ��v�Ἑ��g��ѷ�=�����Ӟ��Q��1~"W���_Ks�o
vҊڻ`وr� ˽����>b9���po���[�{P� �n<~ó�����c4�j7��MB���o���a�"ֺ,>vgw���g�-�o$כ����.��[DMd�x�O�_��g�ݖÊos#���m���<����f�w<C�xg�r�s������ ^?-�x�6W�����z���/��Ygvv>�#lyj1��bp��|��<q�3�����hw{y��� �f��/�1g��A�`�|A�0<�o��8�9SVL�	3ĥ�a��	Ɠ~�&H�gpm?=:w�wA��Ҧt_/�דܾ|(�?n^}��vYn�����^ߓ�˚��g Bp6�uy4]b�@�~9 /X�IF�tG���!%b&1���m�&vU�	;�{��ᡎ�x$oI�pa�r��٣'�[��7��g���o��r�7�V�%�8ꈃ�r`�z@��Tk�w���
����o������"z�H�]�V��s��,��G�lM���N���v�;���`��u"MR�6�<x(+w��������f'�:������n.5�t��{�!���Þ;�N�x_���~ؔ���O�}�؊Yc�G�j�ۍ�q�H��a�ǜt6М�qr��.c�s�ɇc[rvKq�x�-Q�S�v���v��y{Ydu�����7���<hN�P�^8���]ku�m����c'[v��1к���^֚��9�9x�^�M�n�O��/j��ۅ�l��s���Y�Gl8�r����vw9]�������g����ON��%veR��#�R�UX��",�R66ƋDj6ض�U��������N���=i��SfYk�Ҋm;�&�]��������n������F��*��H4�p�4�w����R�`�~��31��P�KyA���H��L��j�mc\z+� &��z*�B��U4��׾�8@�/��2F[�9N4�<o�{�������[��]�$x�K������%�!���E�|^�>��=����T�}�{���Z�ޖ��qSLS��*��� 5Ǣ�,��UR�������>���AE�(�M�,�mX���ŵ��'[q�����lݓ��Y㫢q
LQ����eb��)f�wk������v�UM-�)2�&�)��0YQN�l�+���{[�[5�FsR��uD~@����[=�~� �����TE����Q]v���'�6����uш8��?sV<p������dQ4"�TcZ�TX�h��R���BE�R����W���zn��>�N��0�-��l������B�(��U>�}o%q�Kz}T�t@�����d�
�� ���eZ��2�,�����ž�n�r���C	�("����Ƹ�S�����軵w�U�;���s_�����2�%�	��<�WI/[�F��yb=�z{c^��M6h�2h%&�2S^�ޏ<�z����=½����5Ǣ�-�@�%�Rb��-ޅ^��*�g{�.�i�R�`�\��Ƕ�Ĥ�m���)ҍ��TҶ�P���d�bo�0�7V���#s�:v�|�Ԅ뿆��f��l�`g]�W������b���7ƪ�}�����\ >�� �mF�kBF�Q�U6��`�ߟ_6�U(^΅SJ,n��DAM���7u~���	,�S&�=B����w���枆�a4��BLӥ��U� ���Sy�����K� ��GI�BF1u�FGk�GFB���q[�P��]��AƤ��bP�M�q��m0X��J���z�����O��]�y��� �*��H4�q5{�3����s���g�{���
a"��I�С������>��ދ��������ڄ�$�E8&���<�+s��g�<�������LFD�z(\�L��ջ��{�fW7[���e\�e��e�Ф͉����=��3\���}	���9=�U}��Ą��Ƣ�E�U�^Jڈ�V�h*��j,IE XAd=�w�`�k9�>�AI�8�jHT�����T���̬Q��r�`�wv����7I(A��8�b��Ӷ����rݤ��p��q����C��9����0X)�1�w�U귆{��K{���32amt*�����l�ʎ�&2�����޻�y'�v9���ޡN�fp���
���ŦXM�E4e��w�L�8w�U��>��x�U��L�U��e�m�m��K��� =]��F�TҶ�P�]��>�
�Y�� �p��(�yx�{�[���@�S���s���}B�.ǃ����}�>������f����s��w�bݓx
z����C�NHu��0'�n��ɘ��������$�1���Xqe�	=����.��;�/Z��ظ�]�������~��n5�zв
�W����.Ez���G<�qƹ��b;�j��tn�\��8���حz��c�n�6n�ў��6�<v���=����vnN�Y�s���`;N^x;+Zd,���e7��秸�[y�B��rY�v�ܻ��k7��,c�=���7��Y�nk%>r�HD�=���<�s���kŶ5��b�Z�X�ڍ�-��ߞ����������q��v�f�����c;by#9���ݻ8yS��Ѻ�U�-m��^%8�W~��������)�ޑ3*^�|* ��'���̛]�:!�8DBpD��S���s�| �zz��F�TҶ��W �Ѿ�(x@Y�����O/���v�U\����r��wv�� �ȦmA�1N�>�����q�K}"f}��2�4��g��Ćܑ��8�oY��7-��{����}B�(�uT��Ù�r�b��q�g�q��z���j��z�¨�]���ʩ�a��læ�.\9u�/�w�L���4��Y��+�+k��r���p��L �����}B�z%綫������_y�s���Ⱦ�=�P���YWUT"T�n"_!���j󴭞�6y>Q2{[�銾�sM��.2w��:,9�r{���m���3v� >��Qb�b�FԑB��~H�~>���8|rc��/«2�!�bH�h�bH�O/<��z�'A����uK��:^9�-�E1�ʋv��;��ُ��wl��'�� �?yfM�w�yD6a��l"�:K{�����bޱn�v��M+/cb�.�P�{�9P7#	�p&�T�a�H5���M�R�&ػXs����u�N5�Rj�㝵�j
��ox��W��S����L���L�Y�p�`�� ���aI�����Uo'��|re���7q��|��� ��xG��a�BP[WR}�2Nn�(>�>6={o��C�q����%���a��u���[|�|_F����F��/b$p�K6�č�зGd�"�hйk��o�����˭Uo;�8�"�� ��BEE������{��u�c��NfHbq��m�g���`�G��55z}ʪ}��{|*���E�	���KAU��Tׇ����;���9�"mxU}�z+
��Є�Ӥ"	�����^3�v:�8�mz8������.�k�=���p�L��q��T��2Nn�����E约��xD"��i\"�5UkOEh��
��X��7����ڪ��[�����4�&7�x<�g~�_E}n3��&�w���D�@P�e&*� ^���9��T���i����{O�l�'�Jݞ��S���&_N;�頥�ĵ�ʨ�g�j���{�+�,�rBEl^�]-�	ӫ����dFY�]Y�<s>��z{�فS�\,WPJ�B,��k�3^�����g����	���Q��q��������zDɥ|�<��@}��a��ؔPI�X���_m��q�ӹ�b	�]o���n��غ��ڮ�㋚!BM5&Mc���7�ɯ߶����Fw�k��k��`��`���N��P� ۇ��]ռ��+���3� &��!�i��%�,���i��S����>��X�k��T�^���P�6�A�S*��}�y��Y�j5�D�K7B�� �{�[�ރ��H��pZm$ٻ�Z{�S���*�B��U4�y]ͨ�9Y�� ������-{�N�k�=�d���e����f���}H�j�9嫝�I|+��7錫���	Sf6�\.�&4+�m��p9��a�B.�\�y�n�`�mP]+����C�7`{�oc.�7��#��9�4�܇0��*f��h;�T��_�����x�k��Nnv:�'L0�5<�m�+�N������ɋ+�]F9��&�nOlO��[#���'u�p;�"9j�D�h�
O;�]ݬ{*k0�-�n���^wL�8�v�؍��YE�z�����׈#N�;��_�F�"�4X�m�m�ۻ۷�v�嗥�h����=x�/]a��ӮA]'v֗��e6�]�u�v���Bj!�4�p�pR/�]����gv�:Q{�����|}��/{���4�L�v�n�*��
����Ɍ���z�LN�}�l�A�`�ت1��54p�����Tʅ���i{<#�@(��0�8@��������)n�*�V}�)�����eZ��E��Ma���fș���l+�Z{ʪiE�r�EW����8�1����`��J ��:��<��y����귧g�S�n{��UyJ�b���.	%��ŧޡN�no+�����������o{��8Ӡ �#���=�U�U�Ě�}��������Uʣ�_��˼��o�1�6GoJ�vi�}�2 �|p����]�n�c����ۉԄ@b�{ϧ�ʺ�$�hA*"1AH��k�uy�}��Z��߰gE{9��1����m����O��fș�S����ii�*������h����3�URw�{�����F��]��|)���KF�A"G���L]څ�Ъix}��]ͨ�.R���c� >���Q���0$�Q�[5����'��G6��Ɠ�x}=��5E�rܥ���sL8�!I�v������]�);����.�ޅ2o�q�
i�%"�������89{�ʪ���*Tfg+��}x�g�0�1��qq���`��y9�\ܯ���͢^���B��,n���o,��<cӲ�|�j�;��6vS�א�*��L��o#rg���I�4 KG<���y�8���yv,:O
��Ll�B�s��f��{����XzƎ^9����?x(�w-yl�3����C�ʾ�C�y�00py^����_�~�5io��g�l����
�FB�PzX8qm^U!�db)�fb��mhBN�˷�[P$u��U��ʳ��;!��ẹ��IF��yb���G�ș�%ɝ�'�.�.Vſ�1s�3Iw�����A�j�|ϺB'v7]+f�Ɂ��nա�#T�O�FD��F�� ��J0B�<v����{�Dn�Ct���n��"��s�]2Ի��A�zn{e^�M��+���\��9'n�Й-Ě�ѝ���aO�I$����eԽ�A���/��!ˉ;ۛ᭷�����ӑ�8�7�IX�>�N�ugGu�ҼQa5�KڑLZ{ca��k�MV�O�ګ�Q6����38�H*�����F�g*�<�®���M��ӊc"pT�
�i��rrs��gj>�����T�G��@���<�*��و����{�e������S}�ѐg�xY���2iu3��sn�2�#	f;�V�m�Ź��=zn,��똖��"D]%=p'�ͼ��F��pvoj�K͉��;�N/�.�Jg���xiʒ#�ȧ��f�����n�^� �r͗m�'5?>�s��yd��X�=����<�u�*X��٫�,��5:��\c;���<
_׎;�B��`�5�M�H��)<-->6�r�Od��G�	�FK6�z���؞���Sr��龜�pr�\���l�F����=��.9OJ���޸��,T�c9z����۷���;�F7	��K7 �$�c�ذ*Nw,~ӎb��4V!;�\��P�sA�|dMm8����9�Ёw�۸��{� ��چ}^v(��NzHE������8���R7��Ez�ټ�^�1o�B��nU�e�G��K��x2i@�0:ʓw0�j���֝�X����Fŕ���kM?]^��	�\��{Nh�釸nxs��]d˹�-��\�l���A�!6F2�?XNu[�^S���F��ҟpP���K�@R)?z�"/ZI`od���K}Wӳj�
Y_�;Wr��i\=F���8AC7Z�,k��'ʓ�Cf����lX�7K>K��6��K�m���᚟��QCNui��&����7s�\wݯ�3��+��(-�{�^���pM��pi�s�bAQ$�yNž��ǚ�1�}>2��R���(�>Y�OK�/�{s�.�0ݴ��Eء��߸-�y�;]{���d�-���z%�[�����%���t3�ͬ�����78��֋��g-�5J_!8�����G@��1�s�nq����NK�*�g�3btҢƭ�}Z�W�n�U�A��*���w�s���V(���D�+�V6���W��X��;ӧF���J�{{����pfG������;�;7�U<�����>I-E"LHRpji#�.W|>�U*�{�Ww}:���ɴ ]������N$`��1h�G�8�nM�7�������E}w5ө�N�BE5��(��fV7�>���.�J��Nl�e��誚m��mCM$�"�$+Wm��_��fd��N�wu��͞S�C=T/yw�X�l �&\)1�m�Oz�[g�Q�������U7��ww9z�j���}T-{��Ŗ����UKN�S���np˞��7��O�]�SUƍ>��]MwPP-�U����3U����ysc{~��f~�����Q�f���f���9�V^�:�m��DT�D��$o~+ۏ��7�Cr#02,�76�.J���Y��OW��n���nl���;�23D�``�5��k�����w�L/I���{oMru&�]��,�!�	6��l�y���*�8y�
��| W3��R�q����-�E�0a��Xv}��m���,�ť��T���z�m��ރ�hd����{umQ���h���*�ly]R���]�<��1�B1�T-�;�PNN��ߣ�&Z������4�}E�Y�$pf#@�D� ׺������T9�wǙ�=��Ji+[�m�����$��I�j�c=��d�
H��&Vr���w�Λ�7���fw-�Q=r/����os]]����dNѦ���n���6x�$M'���6,��A�\2# �H����u\.sZ9��y�u
dA��y֋؊���qF5ru��׷�dp�����e�p%a��nK���R]{���Ҡl���u]�3�^T�n��s�W#���9���vp;u�{m<��ݛq;N��3��i{\�Ɗ:� {瞵1�xn�R�}\X.Ѷz�s�+�"�.ܷi-�ba�l+����u����/^�<�zz�;�y�xO��Ff"��{���ŷuO�����m��g�h[���j�"&8v;kӒ�]�����%Ӌ'J���s���+����SMڝ� -���>{��ϼ~�B��r��{���~����f�r���ߏ�U:p�6� ��p���I����/ͷ�|"�Sw���� 2t��3&�{��j��;:R�j8�qq������vd3�^�lk˸��]�gAי���"H�Q�A.��xv�s������+�>�7gWpfL��Aw���@��j�K7G�n�k��E�v,u��r��Kv�=�{V��7g) �*e�Pm$�fV4|}F���:"�Sw����ٙ����w6�1��n$�ZL��V���S�E��3�N?X�N�s7_Y��.�ꂃ�֔�v��rn6*�i�}�s�|p-*�����WA��۽t����C
�M�Y��F^��g �q�k\�+�mY"ȤY=�sB�Ӈ�Ю��>=F���U�������I�)���Wm�x����k��| 1�,YVީ���v�s��)ZL]��I���V��>�sm��T��>g7���{=�l��	�	��m���~>��ŕ�� k�x�y�|�b�ۇ�u=���:ǽ�����qE	Q6��V��m�u��ʜ�mc���G\���V�-m�rF`�YiK#	��'��T���Ү��j��H������um�zbц���$�q"������ɉ��W������od����UM�?w��MHB.	�ʻ�zz�s}�Ҫ�XɄ���񨛎8�׊BJ���V�7����-�֟g�7��:V��X��GN�~��u�`�ܙ����*�iŸH,�R<Z���DDY"{�ֵ��y�;�1���Y0�bM��o��~>�r�{ª�+�*��|.�OyuDf8�IJ*ܓ^���}�7g��M ��ec�����5Ǭ��~ u�x>��\�T���ci.xT+m�$ҳp�ɍ��</\F�=Wb���tk&ͺS_���o{�]ݼ;B��ӓ�ׇ�e�ϔ��[��}�)�����P���͆s�@^N����oW�R�n�J��}���$�E!p����7f�.ߦ�͓���6z���`˫p��U�[��%G	&ڂPEf���g_�ڪo7���xv�S���Q=��&�L�����ՐB�cL�{2��s�P��V¨��I�OJ�P;e�I�ؾ���s��̿]���_��~���Q([z��������%�ZMBp�"�ی�wV�� ���̬z׏�ܥ�©fOC��yL�DL��.D E�BTi��I�N8��vY.���8�D�<]sg$݋9�T\I�b	h��ǧ�U:q�:�][~S�G������X��p�=6�D��(6�e]ռk�Y��dΪ��UM��Wwo���U^��p�0�,�R6≸��5�)���v��X���LOw�fU�k��n�H�z
�ь�ۅ6��P����2ޞ�T���ҳu|>>u�����x6	�\�&cQ������yx�(vy{2qi~*R�Ҫ�mp���S�dJj���d�]]z��WR�v��Y����s����V"���շ::^��˕����,�"�����~���{��AZnm��H7U���X8wV�QW&����yb]n���t#��nڛb�x��i��9�'�v�Z��!�
՞6n�tP��p�:+�ܳW3�nw��=]��z�8[��<�N#�\��s��p�K���Չs�[e���7�yS����C�v�	���a�衺��`�v=ki����R�+'�NP�8�\��ٻ�ןh��dax�z�ߝ���ˎ �r�l��T��Y�b�i�u˶2@��3֘��Ѧ�6g:�\�%w�ҍ�ߕ�Z����J���1��2���z�[��
��IB�&]��o���ޏ�2�{�]ݾ=^�t���]�}���^"�	8I�E�)����]څ�Ъ}��[�^>Óm��T��tapXe.$����
�5@���<�l>����>wޡ�g}T���r�w�;dd��2RI»�x��sm����-]����wa糧w6z��Yģ����ph	j�t����ډ�g-��F��M�ɥ�]h6�$c����M��������6m�=�.��=ޅ�>�y[+��rm�{����Re"�E�(;Wm��+Ϝ'��[j|C��_m]q��n�%�e����е>��ܴ�����݈�|7{�1#M�ྡ�V�ۣ"�;ٞl�T71�������:�UDQ"�q�e�Z۽�n=�J�շ�{��}��07�	�Q��6�,BL]͸}ޅwV�=f���gW���۟}��wa�q�	�Ѩ�;���O�ְ�[|��"����b�o���w�fU��Tx���Eٹ��p�UO�;�31���un;z���o�}��~û��?��X����õ�&�7u���̇)�pIۮ�X��\)�Bbi	C�y�=�SNf»�o%���������v�����!�1�0�/w6N�W�\�oZ�um�G��ێ�����'#��m��m0�6�p��޵��76�.J�'UU�K��3�@��2!�3�%��G9E�/�����q�+?8��CI�˪��V1X�*vU]E�ή]�w_gu�I�s��pɡ0X��h�D��{<^��>�:wsa�l�0�,�R6���no�wٞ><����3/!���������s��\��x_�
�F�p8m�B�v��E����}~����R���>w�ӳvx ����i&aBc���.K7����M���	���j�Y�f��b�<�!��%ApZcc���Uuo��nvN>��Ulݹ��/wv}}��S��Y��	��qwV㷩Y����>�E:Z}�@�l/W����P�!�2�aa2���z�*�Sy�U�����`̫q�z��͓�N�^�[��$&6��f�P����2m���+���q�77U�=&�c�����D�Vq���7�.�zk(�
lY��l��v]>��F�G�IF*��"��ZM �*㽨��B"m�Tr��Ш��9\�f��o}���uϰ^QQ�#	 (z��sd>���PDԄ��HEwV�:�T�� +�=�wov����T��:>1"�0��T���'qh��[�[�+�Fҝy���.uu�u�:�fa��JI8Y��Z����o
�T�p|�U\�9g�`̼���� Bh��H���[x�c�~}9����w*�w�]�ĸ� &���H���XPZ�صv���U,ΡU��㻩Y�Ktz���͢I����I���|���,ʷ�x��ͷ�xE*� ��噖�g�W�n""!-���{�z�6OUٞ><����X��p�z�[�ZZ�����85m��ɸ�26��k^�r�
ݼ�H�q7�X��-<�;b�`�nf"�YlR�u�O~o{5>�&ؖS`��{�Y�oo���1�ä�����E��ͨ]*r4��@7�Up��hlT�6U��M=�ڢ]/��6�tڱ�wxb�z�K���1;t �b"�b�N�7u�F�N��/
�jz������=��{3}O�m�"���s�;�.w��xq��Xb,�.D��p�z ���۬G!.�2j��&��RS�� �Ow��ᛨz�h<f��9��):)�LT�(�T�=�$�7N#FVТ�����ߵ�ɳ�qԃ�Z�{b �8�i��M�we��v8W�Ed��E(;4�b.;!�D\
�ԧ`�ß�[��|oP�ܞ���0n�֟��ʙ(�\f�g�i=��F�t���|??h��<�z�:ވ�j M��s�蹥o��_]����D ;W��ǹ�rq�ԏ`�SM7�P7N"Vi��ùm�v��f"L��z½�d`��/-�C�f��N���h��r�}��{ђr�Gv:by٠��\��[苤��y{Rő�(��!gT�����>P�p��6̝�{=������`�q}8sC�/ ����趞���1�{?y�_{��m��-��H̙��95A7S��5�ok+"]`P1i�2��ʀ���5�^z}�n��=7>�T;����7���h^\�L{�����})뻠�&!�*A�p=X�P�)��C4�fN�i��ܬ�'�c�$<TFc�����������9;�S{��3x��Ѳ����-�)L��q�g<���Q��nqǛE��h%��b���f�n�]��u�tA���Qh����km�݃Gl��ls�1��q���'G>�qd�ܸ��E�n�Bf�s��G7'��g�{bw]f;H�m�Wa@�]���N�m���g�dp���-��!����sǞh�oU����c�5�k�����On�<]�{w&���g��6�·��;[s��+�����a	$8]:��Y���X3�1�\�n.�)� Me�5pۜ�$��n��p󎕦\'�������n�Y����=��C�0@Y:�+�v;;=n�\��Ɗ-v9�l�nn�[�{cۭ�{`r������ݮp��4�1Q���jF�X�-�+�%Ş�
�\f���b���c&͘���חr��8;`{LvM�ƹ�z�Rǿ���֙V���;�C�����\l;�]�������!7=�|B���ܼ�ö�=�^[�����t�N��*��F$�<=�[�o8{X5\�v
=ZCF%ŷ��ݘ��6๥ۭطj7Q�p:��q�VK���ݳ2��:e����k��kE�l�:�0���4n��S�,ˆ.�NWZ)ns�.Fy+'���Bۏ��1���>��t�u�����ݬq�������u� Z����cg�Zc��=�k�^ľN�\�p�7�����!w������r�Y�p��n��-�Z,x|γ�<�F��#��(v��<�����q�|v�pu�ى�}����]S�3����A�g��U���w[n'��].����R�����6̧[��.�V{c���������in-�{s��;p�n]�z:�6�ڲ����vjN�vy�[�0콉w\j�v�kK��Xl�]�v��p[�����v�)���-ɹS;<�Fm٪׸�Vv�����a��Q�c&���k<��Q/x�qS�NTSP��ԋ;�����\�f�W ����è��簧A���9��jv�>w]V)���D�v��$�2 ba@�(�����o�`Cqw��USݳ�H���H�L+_JK5oG�dh !�P�������}"��n�'��r\��Q�y�<W;�c�i�q�ɰ����N{���m·sC��C����3޹��	�gH �h���4A){��7u+�5e�v���tnh�YBsI��p��cQT��XɄ�QVp溝�����yH�o����A]Yv5���',7*rqݍ�2 ~��d����G~�W�v{�L����q�XG�@��iKM�Im{Ҝ��"@��A؅�|8�`�۠k~�qu�7贑�4��M
2;��lWV� N��-��L"����F�F�=XP�^�c����v��ň
�#"�LV�P1,�!1A��u-�W�g=�	��߅Fr�;}(�k61�ƙ�%5�L\��������?���'����ƕ�[��LO-���r4�����x�Y)�=��6�d;h�sVf�o>�M�#b����z��eg�Q�!�7D�(A�1%{q������-US�q&4VY P�"bɺ�#]��$QH�c�Z���؅fO�X��F�jlу���i���8`v�˭ ��w��^�kI�"�sM�,��q2Ǽh�Y����?=��nv%�F1�+ �֐����L��������шa�Gc����N(��,1㾹{��
4d#;}�j�3oѷ��s���fB��Xe����PFA>|q�2ӭs����gf�]v.ی�u�U���뒯L{�a�ۋ�3����т�u��W��Lsƻ<���hupEʊF�{Og��V�`��q��u�;q����f}��z�Wm4nl�y�ݎc��fm���Ë�᧷+ۖ�e��p��̚1�k(quw���Y;{u���앰g����.���6�m��{{���"�����(�d0F���z=��[��^=[Ӭg2�kS��;c=:�|�e#�Mc�qt9kW%�莮�ɗ��m�)�������g���}�̼����V�Ȼ}o�Ғ(�1�!�f���X��VLOw�]յ���nm�S�+�|��OGA�����{����h�͇��=[���]�珏&��{�7oa�==d��D��Fm�
���%���Ij�
UK0j���|�}�������(I�)�Ye6��%�z:�����{d����sc����P�N�^��L�dS5�r�����n��rA������٬ܲ豗���* �����i!�[���wv��X�����=_�9���ߏ������`I8�P\���p�z�׷p.�ho�WR����4�}Ъ��U�l����r"����h��ݮN���}?HuRNx��1�)��{ �0xmp/Ǘ����xot�OkY0�Q �7kY���O�T�`�~ f=�����MCd��a������Q�H�GS�]�w`˻p��
���	e����	�5m�B(Z�g�י'�����}b�o���޵�*��~![pJpR�#[�y�b������B̬kW��m�w�q�OP���1	�C&(L���%�r=�o^�ǵX�B��L�\j�V��[%�[E���AfV==�sn;���͑N��UV���ѻ�;�Y�Ċ12a$�+���w;�� VL�;��Wm�=�������Ug/���@���QMa����z)�;ݱwz#zEٟl�ɟ���=�z�lk���A�y2n7�˓|��
Ƶ��=������¦�%��Xc��M_U�w!D�dW3G����u�o�c������Ab����y�2��:޷Y�y�ۻ�W9��$g!)@��� :��T�t�����hS���wW��̿G���"4�Q�mC��P��M/�;�]ͫ�u�-Zt��c�UO��>��L��,��)4���K�
u뮗�ݎ7�K�;>�\랣r֊)�妅�"1�5���{�������=@̅�������ǣA���ʓv���\"����L�G�����X��q�Ԭ߀�d�r^f
%��aū��B����Ю�c���ɦ�]p�Wm�p�U���J�s|�����>��麶�ƝVE^+����'�U./��a�c��p���^�Q� �C�hb���&�30���W���Ov�p��t�V��+��c�Ux��L	���F�o%:�����5�h�(���h�z��6q_�=d�
d� h�܁���cޫ��n��f�Ř��y]ݼ=�w{�U�x4�b	Ȕ`�bQl]NӤ�m@'��U�����n�K�mHk�ny��e�Sj��X�x�R��wn{����ɏzj*i�\)p���L�I��]���ye�����.�nc��Y����<E�3��<#��FʉG�h}�UJ����>���|/��{��UK3�[-��2%R	ݛ����V�|��T�^틺������fU��R&A�[D&��M;76�k�v�߾�	ޏ,�ǧ�*�8��Vn���7۽qԽUh��I[��/�����}Wսà��PԽu�ia�2�o�V�ݍ��̘`Kz�f��3Φ4�^��02���?O|��~����+�\�]wg�z��h��ڭ�����kn���/5�֮��NK�S	�൑泷^ӻu���gB��˗-��se�ۓ`����k)�]�����;���c���u���˛ca�wKІ��O�Kb���n5�Q��z��n�]ɦ�T�Ge8��a6���7fwv�����6����ru=c��^y�;�ם�ϯ6#Th�E�P�����_Wnͺ��Z��2�<E�<\Gom����܊�u���m��^F�aj��^�� �/���߬]ոy��[�����ɝ��v��ox�%��I�"�#]ռ=�.��²c���7V�c�i���w`�����	�Z�LI�	&»�z}>�sm��� �2gz<����z�۷�9�1	���A�SVn���&u���̝>��̘���̫� �^�aɶ���H����-D�Z�o69]ݿ| �?`�y��z�6N;�ٻ=B�p΄�"
�4���hzW��ͯ�����:���#�K1�8�	i&�D"@[���g������sm���d�������e��Tfpn͇��=[�����,rw~�j�����਎�y���]v�A�O�B��7)K���vOE�rWi�����Z8���ȋ�f�*�IG
���zk���s�i��	`���XЖ�5&�h�wF�2c3b,#����������n���X��p�+�������D'	��BS�sm�:��Wm��+���d���f;q�z���l��\�Zm��!�n��}:���n��]ռ==f���� UoVxF��Ǽ=\3���.��}��]�~ }�ZÕ���wou�������<���p��"�'5b�lg������vS�[���R�-�+�;WG6�i6ͭ>�x��y��E���G/}T9�r�����g�̗!e8�rEN5Fi+X7���'3cޱU+���]��Ϩ� &�����d�Re��m�n�w*�W��+��y۹���n˕��o/\��� �w`v�"1cG��5�ڌ}��*���C��D����z)���\f Wv�;��6�w�pE^73� �e�����Ž*J�1�1��)Ƙ�E`Qb�*��"���Z�s;�Wo:y�!��i�.LUO��Ｓ-i��IZ��w~ ���ݬ~��i�ۆ�`�ᤘ���*��^����c����3-�9޽�~��֛�$��d�!�.��h̀�}��>;��7�{wp���ⱺ(����)HYj i�4�o��{f���M�u|>�c�{Ҩ�%��$%�S��n!$B�w��B� �����Wv���P�+Y�~�9�{�Y�M'�Q5UK7ޱwj;�U��l�R����R���!@�E�A�#��P�>~�i��-�����9UWq�,귋���\:z���8�$�3n�=4�vY$�<��ɷ���Nӽ,��Fw�^�nؓ�t����uo����/'1���ou_��a�AdJ$ �	�ݓ1b�!uԲd�*L�����+-n�9!0�$�� �)�3I�S>��_}�v���y=�|]��߅P��|'������Ң�Du����m�Hv�ۋa!{M�-�u����`��_�]�ʪ��u��Q�Ҩ��[g��N��y��G�BL]͸y�*���y:}�ȹ��uxE���G+��̘ް����I'��>������VO 6�v��{�]ո��� � �An���>g]w��v�p򻵙�b�����{Ԭ�$w�/3�d�DE�����������Y��O��nm�S����V�9�]g.��9f`�a�=�V"���Eo})��IAGb��tf��)��,K:n��+�|�V��|Ǘ�3r8��n=�W�]Y�3����V����v\���Ƨ��V����t��[��N������;%��T�3�(Ó�epAv	�י/CN<�s��Ӎt�1笛���yX�<��c���q�bMخN۞}���Em�� �"�m����۶���#�k��P�y��n69Ӝvkek�9.;X���󳻆۳����8m�|T�v�ӹ���a��!s5t.�[���d�Xc�7p��w�=]���H�d&bO���҈���R02@�$ IETE5�+��j�&r`�hj��SOn�����hc��v�xB:]i�%�9%0��.A)����un;����l��?| ���=�.�ߌ�(�l2����e]յ��Y�P ���]�m��ޏ=��y��Ux���|�rS���%4��um��"�S��b�x|LN��̫kW����x��p��%�d6�lw~�請���ێ�SN7v����Uw���M���� �`�8�*snowV�������98ީ�n�|z�wfרR5_��?�4�� `0̽\>K��=�n����i�ͪx����6���Ůj��M�D Kq�;�\~�54ݩ�#�9��/��y�U�[ޓ��0K��D0�M;76�)�΍�L$3}�39�;oy��}W7<�^��#�մV��`�B�H�r�SN��;F��J�ګ�7UYU#;5��;B�r�s�7�T}��hA�(C4�&���!'�]fw]�dE2,��F́4dA4I Ѣ#˽���ϗ}�v���z��[˿{֐o���rAm�ٻ>^����7���}�G�eN�/iٶ�Oxwn3��0�i��je]��|'˽�2mǻԬ�[x�x�w~��}�t���`�p�q=������od�U�w���o{�]ݾ;�.�߇�>��C0�s�
��Y��ೈ���)�4GU�nNu�+��mQ�<]\�^M���~~��~�n��u���7�� f^>�K�'���	IDTp-�o�u?Pwg��빷�R�um��/�}��L	��Z!��$��[������ˬ���g��]^���o�Aԑg��398��:�ww��q]��}��-@�*�^�v7��'.#o�kyH��[*1fu�L�A��d���wN�]�q�u�I5��F��o7��eG)��=_�������{_0F��;{��4D��9,�s�ϴ�E�}�I������Z��]ԃ�+N��!VP�j�M����d����x31� ��`Tn�;k��q7���-mVY�*Ȇ7�G���װ�̃¿{H���|^ض]xڕ�l���{;���+�#�q�5	�?e��L��$b��L`�֗\b�ܵ#5Un�R�i���F�����H������Wꫢt���p��v˾������m��T@\^�j�1�]Ƚut�^Io��\�{/���'Y��8+�h��]4f���
�g�w��%�ԇ�}������r�++}縵�����~�O"XTu�O1qb�N�Y{��!{c��}7$�/��y$��B�����:�b��M^��?~>����Z��lS"�U\�U�wfw%w&#��$0M*Ww�����U�7ۛ,<�3/w���b���"���«�D�G����\��L]���py����{��;��8��#�×��)�p3�n��-Sg U>����Z ���ca���.{+f�<tm�o��[y�=����?Or=r`�q@@Cb���Qf�(���mh��2%�;o��6 DU[/V^���f�m@�u��h��3Z���~�<���{��Z����~
%#�׎�6�30
m�3��3�'���{o��л�xA0c�m���:����RS�#�������xk�	�!Zǉ'D�d����JU�v�B��]mN�{�;��k�h]�D����i���1�I���T����g���R.�^�K�#I��,��sA�gFT���8.)ر�q=��O������?��-H�D�xL����|᣼��À�L�&��P�h� }3[ݱk8�^ig~[��9��~OO��y�mئ�����~�^�x��5Np]E�憚H�eB<z�ax�L�F���c/۴���L�)kA��f9���L��N���N"��M�w�B�4�M߼�WD4�Ci]��_��(Vr���)��:骊^� ߊq<�Tf��0`[�&u��ct����5�a��"�ch�y)��P�q�,��$��"yh�B��@a�0�+
�B5�Vȍ`�# ����Z�Yw`��P�0��V ��C�A����
;�x��ް�Zr{�'���/$/A�or.���֤���v�gf�	wFȰrc9k�����<l�"P���QA�j�E�b;`�3:�"2}�� gvk���n{��_��`�`Rh�th��c�	��]�e����M�sMQ�
X�)r����I�t��n� c�ʾb#���T�[��F8d�(�ཷ��[$�����\7�?9�h �B8N�
o�<��ٚ�`íxf�v ��s�T����XIuo�����,��9rk*�r���*(�"DI1�ґ�E�Q��!D9�4#G�9Vp�wm�qWwn3h.l�np˂ �.���ހ%޵�*��=�-ݼ��-_��|�l=��L-��
�I;76�-�v�߇�mw���~=�sn;{�V���U�y�@��t�"P��;v)i:^���q8Z. Q�6��l�h�-�������.��<�*\�χ�edή��̞��(�R���e��Wuoǽb���&=޵����=�-ݼ�~����]
�6���)��-�wV֯/Y���o������K.����^��΋�%�YN"��G����
���w��v�ޱwv���Wunx��r�^�'Q�����$h�p���{�Ps�v����4oA,���һ�X�TA�w>�*��k�9�f� �I&���$$
B$�J!��~w	��0H����0��{?k��w=Ӟ�J�L�L�j���%wv��×{d�w�Y���N��߇�o��B1��p�͑ݼ�{:�u����r�/9{J �獮��u&7�@� �"��S23�g$��Owm�\���\�.� �w;=�]ݽ��-4�d%�Zb�m�oR�~�y3��=����wm��W~��;޸FB�XiCBA&��o��]���y]߇�d��`̛q��+7V�wI!+q6�A�I-��|�љ������k.�s~Bｿq��������G
J"�{��Ou��������k2�q}�t�����A:7cw�ѕRf��\�3�X�R��m5i��g�@�x쬰��ܨ�5�[
���
�R�&��yg�W\���wl'I���N���7�4JvnE&bI�I�=/#=��n�`�������VI�-�������c��Gk&�VϠ�q��[�gr���o������9�����hÉ��V�Y�\k���n9�&��#]�9ZD�n@:^��޲
�:SΐwD���l�+�o<]W(� ��0m���;�����c`�v+���cg�"��e�7V���gE֭l�:�{R^��w�o��cM)����;t���\c;�� ѢI �S,6�%)������}�]0�Ws��O]�<�u�k�e{Vv#�鐆�\뗬CC"pA�����_��76���v������fd���]ͽ��J,&	!��2�j�շ�v:/� '2w�軻o{�]�������U���wJH�Sk{�*����w>��ʏw�iڶ����f�0�uF��@�;������y�����76���v��>v��ff�>��&d0C(�ݽ��w�͏�κ=���wm��v���z=s�`sx�Ny� �X�M�z�\���}�k���u���>�ke�O#����Sӳ����v��N�Wwo�u���edǻ��nl���ߢ)��f���Λ]�_X���&�q�\��'
XG&�?�~}��W:�ם�#f~Q��(u_e�"З�^�!L�kF��ޙ~������=��_�E0EUG~.F0h��s�b���6�eݫkW.�sm�~'9}]�D�.B����=����hݻq�Ԭ�{��ɞU���v��軻|gD(��P\0Jh�	��� %����oy�]�K7�����u�t����Bm�����濔�������w[��eו���Y��� �	�#
��J�t��s瞻�O^�#ɵq��m��ЋȽ��kb"���0��Re��M�1��wv��X��q�Ԭ��y3�z=����.	f0�e����um��w� y/W�������v�o~��fN׼�	m4�#�ػ�q��+7Vީ��~kh9��r�Q�핇tJhN��בԄ��ޕ5���`�"j��j����A۬�rJ�\�V�-���@.U�uZ5����O(�,�BaQ@H���Wwm��2���w�jL$Ra��	�iṼ F��t��̬9�)ց�g�֢��v�	S�JM�$\8�7�bc�����q��*����/4�0�wsJg�a�P#$�c�{n�Y�nu���Lu1��m�����ѪJ$6�����F^5*�� ]�.�g8oL�!�i�
.����'�	��w�]�[�*��W���U^���&�p"���M8�f5�|}w��&}��v���e���u���ЂOE)I��}US��=����fJ�*&sz{r"!	�1�Y�=B��m�L��{Q�~�A��^j�w�
9��`���|vIy�y,[]�pi[�'�q�&���U�h�5����n(��\N[���$��"���y��Qt`�j>-0��	�饹�f�߅P?zi���2M��wvtU{;i�#fn�7eMnH�|�\t5��f<�8�i67�u��Tz�ħ5��k�l���_�^�+7V�K��n�:z=��]�[�>wj�w	��J1!-��ӷ�/�3=T/v�7�����
�N3v�����"��[M���"����UX�owk� 2^�y�d�g�*�SÕ����I��MCE]������vd=���nl���ӳw¨}����G�mA�)��$[��qwT�K��xu���x�����*�>�}G�F[�]]�E����ݚ���o�N�9������';P:�T���0+A�NULP4�+g!�d�P�"��j�^�wR�O�C�:��2M⥻���ba�S:5mN�7�����b������e�ᠻn��
x�����v����<r�X�kc��۵��z\8�q�<����\mir�n7�����qcv箻
v����Cq��,��+̵v�`�-�x�lrʾ�vn�u�q�,N;pJ�1�wcN\:�r�V䤆��հ��κAWu������9ܖ�M��o�Uu���%^���DX���m���[�Q�&�D"5D��l�Z�Q��Q˵=�85�4�2����{t�\��G#�6���٩���A.T�0����~������ut]ݸy�W����{�76ޯT/a1��8m6��v�o~ᙓ��N�v�+7V�K�����{$�@�nT4��/&'{�]յ�޹��dή��wm�A��w;�`��.6�(]���{�kU���}��wX����	3��*���I%"Xm�A0�I���y��ڻ~�=�n��r�n�n���͓� ��O�F\Fс��" �ջ/7n��n���S'����6�)�l͸�aJB��a(L�ǘ�ޱwv���Wumb���Ug.����{�����h�d�#Ew7��?`�b���|�}��jfh����;�	;��2�� ����W�q'7h�	���D�֘QG���&��N�^�=�G�Z�u�}9�-�z:n�<�|�Z+o�5�FܮEt�F� H��W9��չ�r�N����F��s���{�ʈ�b8P�8��kZ��76�k�v���2g�T̻ն.ݿxt`���ʈ��M8�no��w�_����z��ۇ��]�� 'Wz�2m���A��R�0�׻'����[���1��R�um���N�����CQa'�GN��\�:�=cIu�kv�jXTx0r�����s[bZ)$K-0��	1�X��x����z�.m������d�32�����a�e���a��ǫ}U[˵~"��߾ѻ���Ow�l�z0'�BmĄ�<�������"ffO����FUJ's/��v�C�& 4{vj���S���� ���hDKr�0��a�p4l���*z�Ι�sD�K32�t��'�x��@q�}�}]�����Hy����*��A$D$�$iq�o�3f�����l��.m�e4�&W~�};�`��p��*��ޫ����	����Wo�P�h�M�a��0	��yˮ�Ӓ� �޵�+�>�\��ۻ�� {�ϜDA�H�Z�5<��K��mF�o/sl �[����B]q���IB!���f
h��efV==�sm��T�����32w��v���2\�&�mHc���nl�w�3�@L��X����Tҳ�B��ߧW��p�I�p�d+Wm�+�����߾&=�ZÙ��@3*�zK0�a��C(]��I�w�̫z{�qsm��T��W��5_@���-�
Q8\1:``�Q)ɫ9�;���>�uU�۝���Ŗ���+'���q�k	ah*c$�'����v�՚ɾX�߾����bL*L�A	h��  ��B6���yݜ���)Ĥ���4�ݛ{�z�6O
�u���wX��p��U�[��C��*�.f9,�����m�z7�1=�e1tZ�ݵ䙁w]W<��I`Z����Y�d�|�*����Wwo|�~�|3'&=�R�um�za(V�-��-$\Wo;�_�fd���U�[�ޫ��oW	��|P�➘�FH�Q�X�3=�n����+� -�[���wX��y�b`�
�d�e]�����^FM���.��y��UxUO�=��
.!eDCF&�x���tUW}�������UTY�s)���?����@@	$��D� �I�����3�g	H��$��@2�HI%$$$��BB	h	�!%�����0�$���H@ _��?��W�5�_����������)���?�����������������������۟���9 $�����)����?�� �I� $�����������z~?3����O��������v���7���O���Sm6Զ�ڛjm���ږ�M�+Tڥk-R֛jmfڕ���Zm���i��j[-�Zm�m�jkM�+M�-�mM��jkk6Զٶ��͵-����Z�ejm�mKl�J����m�j�jj͵-f�kSmM�6Ԫ�ږ�m�ki���fږ�6��jj�j�T�Rږ�U��5���l�M�-i��kVʩ�����Z�i�֦ږ�jm+V�ڛm��R���6��SZ�mMj�j[i���6Ԫ͵-SmM�-�m�ٵe�6�V�ٶ��6ԭM�5��R��jUfڕVm�V�mJ��jj�6Զ�m���mM��U-T�SmSmMj�i�SmJ�5�VmSml�R�ٶ���jmYm�Zm�֛jj�mMm6Զ�mMm�jZ�����j[l�J֛jm�5�kM�-T�R�fڕ[6ԭ�m�[jm���m����jmU�T�m��+j�U6��m��j�j[kJ�֪m�V�mKj�j[l�R�͵6�6ԭe�-��R�6Զ��ki�-��Z��m��j�[mi�*���kmi���jm���͵6�M�5[M�j�m�Ufڛm6Ե�f�m��*�Vm�m�j[fښ�ښ�mMY�-M�6͵-�j[6��m�jm�l��Kl�kSiV�m���SY���mM�mMf�+6��m�l�SSmJ�jV͵-i���6�մ�SkiV�V͵-�6���m��ٶ��6��m�M�-6ԩZ�mR�mJ�jZm�i���jR�6m���fڙZ��)��m��Sfڍ�%ji��m�6ԛjJ��jSmEj��&ړkF֍�բ�Q��զkZMT���h�hڴ�ڭ[�rڭkt�Q���SMj+Rm�6ԛjM�&ڔ�Rm�-Mf�*�i���ٵM�m�?P�����~G� I�7=����J?��� I$���1���UL�<������I 	$��w��������?Q� �I��$ $�~��D�@�I7��� $�h����c�(4g���Q�S+��EI 	$�?_����'�~�� I9?r~���o�~?m��?�>O���0 �I���d��O�k�;�J~��s�~f1����������}���r@I%�w������0t�]>��� I?Y�׌����� 	$��������~�������X���W���o��PVI��Q@� ���\@���;�do���  � 8KG��                 
  u�                  {� ��	@HP���� D(P� H	$  S{�   ��{n<^��W`�A�݃`t��>�:7��v��ö;��c� �Q����_YNo�����.�{�壶{�>��/���F��z��죉ݞ��"�U�   8�@,�|[�����;7��[��,[��W�{��wg!�� >]��}��J�EP	��=n�X�/^��NA��`}nϽ�z�l�kvB	   �*�=y�����=�|�=�z����}��{==Y�q�.ϼã�(B�.O��su�����'���P�a��9t'g��/���`z�;�<���%R=�   �)֗�o��o=��a緧�y����(��;���Û���.@��T!@_q��>' 3�0�v�$��q�n�[��u��3`""�p   nfp:������zh3whu�K��{�w�u�;��l��^��RUQD����>���e���hi��`uÐ-�Gv�}�    �Sb�%�Ɇ��0&�1CS�a%*R�F� &��0 �05<j��)F�014�р&�&�=��$�J� 4      ��HI�U4di�d�&���4bLDjR��MG�hh=M4�=4�H�'�}?Wȃ�D		 Z?!$	 
@��$����~��* �! �_������1,�� ~�! SF��*H��!F��@4�$��KM}A������!H�X��}���
��>�~f��g'�[���?�/�g�7�K�1��Nik.��w��P�1�/
w�g��� �d�+*�
�Ǹ@����o���?kx�έ��n�����OqѼ�7H�4&�b鸁�C1ǃ��z��V]6�Z���A>q�i�[ �A�ض,LuGvV2�P��n@�����V�,PDS�sq�d���)z'�b\4��>�u1bX)���&b�V[{; ����� xK�l���EZ���.d=�X9�(ҲM7��@���݃�л-�5ǈ)�� ��Z��Y�掯:��u�Q�wM�EZ��z�ٔs��r�٦rF���f֮+g-i�D���o_��0]��ɊY���hqe�+�yBB��=�5R7�t�WǱO��h$�2b��ېJh�5w+)���P�d����gE:�׊tT>c��L�L�0�w�Ǆ�{rl@��໰���[x��������,s��N�5,6�H3�)���=�r�Z��4��њ���7�
�6D���%��r/t@�m�ro5\`*��5v-�i6�}N4�.�k;�jR�/�GC��2v�,:u�h���zL��Ɗ�1��NW"Z΀�X�7�^����^�(f�A=�k�us��1J�t����ع� 8�h�X�D媁�Qv�^�RU���ל�2o";E�JP ���ov���D㰘2t�˚3��Փ9k%u�8`��A�p.K@m<�뷞MПM��\�y���d��tQ�r�l��[�������-;�{{
1���'�n֑��ҹ=�ˋ��OFV��]�es'N�YL�њsBջ�`����܄����t`���m�_N��km]�Z
-�OxOn�9j�,\�&�^��t컖�ᛴӼ�Ur(�_�)�rJ�KY
e�M�oNTE:����r��:r��9�N-�8S���`��I�<��Vo������;�s��y­�L������9�;ǹB�H���ǧ����W#���E�iq�grx�Q��ܜL���w�M�J����ݹk9�_Pށ��j�1,W$�q��
�Ӝ�ٹY�?���oN�U�:�8��H�����;�1D:�^�3I821�nPMp�P� o�{f\����������$f�6�����}uvs�����C]Z�B��Mc;���n�kSKǬ����YA�˺,�����	�9�+4�V�9˛]y���2H�P��P��@�t�:r�MJ�{��`�^̙���:{]5�]�Y��C#�v�"��O��F����ekΟS���rv;����ڠ��
�p҆Z@@\�����vv)����T���l11�].8˨-��
X�!"��={�����ɒHz�ka}�BU�Ȱ��p�9#ݻe
ni���f�aL3
���Ir�9�	v`3y�����'(��$���f';��41��;��f�,.�X���C3-J�;��V@�,�`�t�P�)0�n5�hׂ]7Yk(m��{mg�4�F�ɇd�1qK.X'Q;�z^�A�i:)�F�#X�Kǝٱ�w6���Y�v���pl"�܌!��p�7ot���r,:�7vπ�em�:�v>�8c�V��w\9d4%���s�qd�pI��<���	bPA���X��4ZV��(L��׌3�w�/�~OC;q�}�"ag0�6�B<�㣆7��;r��e�ծ��a<�`]iߐ�l�.��}���R��v"G���F�Y4AriQh�I���m����-q���VW{v�98�k�6�^v���h��H�v<�Ѿ��;|w�<�gIxf�n:xNujAvIp����3�?j(���]����ˊ�	��Ɵ[6��B96&z���)i���P�:$k4]�V=�w%�C�ȓ84�׊g,O�w�ajh)�� �o%�u��%�8e�V:��y�盨�3�-�kѹ��L��W���h�HD�Iw�W`i������chX��BH���v󠣳�M��n���)��-�W���Q&�'�r|��x`���K��S��Ь(�������M@�ų������7��Z��n���q}x=޼�;�oJ��B#ra]���4��.v�݁���i��Žx�jɬ���\r��b ͢��6r��Ƥ�����ب�$�\$���z�$�e��灙ʯ�v�S}K�7^^[�q��)؃ܼz����*7M1#]4�^�%x�-����By��-�)����s��'I&�6B\w�����t��;�fF7Cy�ޛ�Q�{��W#���U��,8E�[�շJ�E�� ���/4�I�f�[��{��Ks:S�У�nPq,1滦��a���Ќ�WN�L�@���uQ���tH�w��;Ʉ�9�zT]p����ozت�qgp,t[��6�"��˹���t���4��F��������tb�xt[��x�0SA�3�"�l5�peӅt�jv�ӣ��>��w@���õ�ƹ�R�Yݬ���ۙ_Y�7�+"�R�G��xH��0<
1�њ���ȳ6R��y���Xy�j�K{oW��ițL��р�}gE�&Uծv�_��v��+��z6hzgr���~��-�ȝ�gr/���Oc����Xh�=��B��{��^�!����t2��#�^�X�Ojn�+��sj�t!lPӜ\�H�E�4液�o��ݩ�zLۏ#4�.�}�m�/dѬ��Xe�ygN�t�eXW�Fh�.���\&��#�|�>*�fG k:I'Z6gv�[�M1GN#t�.��,t�taM0s@{�4�Xw%z�=�H���N�]݇��4�.�ߘ�*(1�W3������:nG�.m2v�'c��ݿo�˫A�Fw<�3��Ф���q5�C
^�H�N\��'B��wd"��Y��ĠYʍj͓M��Gv��Rλk��?,�8ַgs�sK���f���r�{3s.���cӣ�ܻ���a��v�>G��5lNɡ(�T�Q���V�+��r�	3�!��wA��s�6^���0k7�.,qr��y.�ݰ�!��+u��f�-)l��f[�pG��[A���P��I�����4xݮ���7Zsfr�-:X1<�k�)!���:� �� �h�{�+s�)-}��l����q�������%��-P�C��J�q9�6�8�ެ�M�;����7�`�U)�h���=��:f��ڹ12^�%Q�=�ޙ4��=˳��+`��Z�s�l��f�ϒ�G6��X����U�H�k1�Ʌbk�v>�Pޥ�.��$���4)J�� )^q�=<U�z�����nX{g:�k�rJ֗�~�9l�U�Gݻb1�"r�Fy�1z�cd���*�;a�ٸ�r�㽓��!(����-�.L�rV�梛�����;N���7齆�ҕ[���C`��>X1��C�i�7�ƭLc+,�/f+�`벛9�� 6<�K�3���n!��SI���8rvP
�7�Q�:�6L������>�F*&���K���W�o=;a[l��:N��ݢ�������T�8�r��N�ʃ��eḼ:��*���0��]^;.N�M�~W�wPr���^�N<Cլ���R���RŎ�҆5��8�R3�n�.<�������q��Hr�k'FJ�scyt�އ�rҮꌅ�Zo��dl�<#S��&[��v�#���d��D0�� ��'q�	+��@�>(��^ 1�2 �&��CI'���^2�����+RҒ�p;Es��ȴT�C��G�*�g��������Ǿ/�2���/��ʪ�j~U{u[u�J�i�m@Ճ��o^�����D��u=r2luvx�����lL�`�ϓS`�n���v�뺔�x�������Lev���D��0¶7N#<���9�uʷ����c\�Fl�3�]��<Vֶ�^U��:I��������nѭyst=�g����p�{�q�mk�7\����EOR��Mۛ/����z�$:��DP=Moe�zr�]�n��n�XI.s�����`�v系]=u�'�ܝ�S�wm�A�VYК�^.㈇���'#z�3�f��q�kn�^��/,.����T�LNs�qלvҨ�Z���9{��b�=]�z�<n6峎M�v�uٴ���5��ݪ�w<)��7b5k������[�&����pn��;y�mح�����6~\���c��bOF^��k\����L��W*��lY�9��NL�9�l�Ѹ��Gt�X��G]��b1e9wV4qr�.�&e�Ƹ{���i�ź���agpT�\��Y����v4���zx�xw\q�n��]8݃���s�����j����k8��m���]��F�˞w6��:Z��P�\�=�#Zy��7]v�m�LN�8���]ٺ�F���!�)ے�Y펶�[,: 3����m!���ǝ��9v_7����Mؠ>�=��[��m\�{ev�p�M؀�oE�wj{XẪ�+�i�[<=m<n��ź�1��X�0꠻mτ��S��Z���7h=Jin��3o�ϗω�+YͰi�b���<��6�T����s''n˞:۫���@Ergm�&v]�������F�1�#=��6���wNc��՛���'6�xre��g]Y������v�g����6����؍v��O=3؎X~>s����מ)���h���(#��˹���v��(%۵�:@�`{o&�)nm�z}����(�i���k۫�62YŜ�WE��M�{fN:�{v�<��tx�kb��zZ{q���j�M�;��\��n�G����{����IG��������8;g�kb�L��l��<oi�).­����<�C�rIӻ6�l��=���:v�=��a�bUy����k��U�ݻ8����ɜm�ŵ���c�තc\\�МAs��n�i۟Oec���3�#���)��<s�4lv��Tx�#�+=�\h3�ӈG1�m�a�pm��nf:���%���L�W�0E�ϳԸ�.�j���Hp<� ^��q�S�d�=�7K������I��ö����ny1�ܸ��	���s����L�l���:޶�8��%��rs���86]r��<�06��n�7|��<��vkm���v�D�z{���Q��z���ۉ�-�2��[��Y�[p/X6��k[uƲg�1�ع�7[i�)�^[4QJg!�����cJk��H]�l�s�p�zܯ5F��zF�Z��͔yb��g�V�K�,<�荇����b�l�7:�$�9��[�������UB��a:0�v�̫�g���E�=r3�bu�$`�vL2\���Q�k�]�^���g�DtqkA�Τ����<r�
�璺zz�9�Q�Wvk���T$j�t�D\�K��@<�;=8�l*�Իn���1��۝��m�kgmp:�M��m�w-�N��m7��.n���e#$n��莇Om&���(��e�՗q���a��\�eŻt�S�9�-[��.�6��w7��;U�vxg�G(tlݞGo=�[n{l򷇍װ[���'���uf��;���$準�yᥱsn�(9�;d�J��rrX�l��;�Fp�n��{]\��QYͧT��<Q��aP
��3Ļ��h]��m ���;�;��^�*�;�;�9��Z:�.4�����m{��u�Wq����tn2��t��A�6c)J�ӱٱ�v���uF�2�)����r*��
2ի�ۧf�x2s�;vu�Nza����\�4/6�M��(���74���wg��!2��61�m������ۄ�n8��m�����h��l��u�b>]�F�xy�I�8z�6��m�]��g�۶�q�����z��m]�:�g���R��3�H�괮���c�2(Pp�w6�J��R1��X��v�ON�Ϊ�݇���,�O����#�v;BF)m��nx+��I1d�s���4�*�:�f�L��mx��K�F�ɸ��9����Ϋ���Cn:��C�&�c��狸���=����v�Pn�Yo��X���wp=qتS��9�;ooQ�lA�q�N�����j�g7	�5!�7,v+�ݞ۳,��i��綧��������=��x+�t[�q���i�e1��^��S،��ݍ����'M��n���=���^Wi�e��
��˙��{Jʐ�Pb��Q�j�ܓ�l���[nwh�ջvlX��筌���:��n�z� �&shs�C܉�+ķm�$mϱ\��p+&�mv����7�c\�b:�ɥ��˸��\]>��r��n�q�譓;wO��s��PJ:�j��[��-���M���=g�ʕ���ɟ!�Z�f�w;��msN�da�l�����y��-��%N]<Y���¦�,��w�� �i��3���'�sѹ��6p;�,`��/�{��e1!k5Ν�s�g�q���j�O<s�P��>;	�zK�e-�$NRl��M�&[��>�c��yv�u��|;����<�����w^�zR�;=]�Ξ�v㛷e�ۑ-��;=�����]�u���N�qAsc60�Lvh��s茒9l�#�p��Օ>���x_� HH�5�Z;� �_���+�/�7���E7�t���4��b*�+���Rmzǎ��k��^X�!�4΃!^�*f��f�3q�7Z3}����{{7�rX�ڶv%��E��T=���=�����R��|���Lz���C��7��I}c�07�A@H �gzv5�c�̦}�͗�^w��e��mg�7|��	��� N,�4jk���v�cĝz���m��{I�t��gۉ��NA���&u%l��=��Ucwu|eǪݞ��6�y�~`�����9��;|}�龆#���ӻ�[�Y��{a���ዖƞ�پ�U�Qw;f���[�柗�B{{���9�`���D�1���{2�a�q�OhPR�t"�$)����d�M�Aj��˻�kg;�/w���#L'�܉^���o{�b)-�Gt���lUޜ͈�R1	Hcܯl�j�T�;���4^,��$���;���G}����|M��< �~/x>�npx���N'<܇�\�]���GK}��~o� �8��ۼ+��Q,S�����޶x-��'�f��?2c��ܗ�h�@�{y�{֤��5�A��}�&���x9��z��$:JDi����% �I�����zW�h^j�o�L��,����ʉ��{Fƒ7�i�w�k}/L�1m�Ɣ���s�Ǘwz�{��$5�Ƶ��V��D�	1Pu#q�Ѧ�:�R�ݢ�i�z���vv{P˛s:*�Ư�/ gص�G����ӗ��j�|�������E��o�؁�H�=���q����ϟ�����#��W^榏R��>�E����Csn�_�L!�m=��b�ɽ#bh�z�cۻ4�zv�hͺ�%ԊKY:}7��
*���%��d�¨YGWj]qY��1=s�W=��nk}g���3;tw��ǎ�^�:���4���8�8�2�d�3����K7�8 �y���.z�KB�=}q��`��jv+�}��s��G�ӹozz�3�;i��A���얁p�!�t���(q��Dk5�Mk\m&D'tb��0"�D��fRmL�b0.�6b;�O��%�ms�Å<u�n�V%��r�L�5�_sx�y�����Ҥց�ahP��uw�S�;�ڤ>�=���;��
�V����y{��w.�+�x�k>�S�L�������^ALquw�)�Ǥb��">!�S��;‷�F@[���]=�}�J�ȼ;�.�-&iʔspl�HcH+Y61�n�&p�!d��ر�4�3�މ�6�N�̚�)�bfxg��]���o�tѡ���1d'�����Ą����V����Je%@r"F�z�c�G�gz�is��[�یpĘZo1�6͈H��.�l(ܱ 3�g�[�if�Wg��Eq�W9�w{q���||�;��޷&m�Ӵ^�eKno.ඝ������.�����`�B�xm�7�oi[��
�|�~"��c��㑠Y~bo)�Y�;�F^}�ϻ�9�}�,���]��W�+u�>V�Hm�o�L�������N�n�4����;x̀P �V8���Ïa��!s����&{庌��H�N�ӝ�mw��;�up�o��.����������y�P{�1b7ҫ5�:y��0$g���RD�96��~�]�b��W8�o��ɫ@�gf=a)��1�)⊴m��e�#4�����}x%���hx�K�b�z���Lރ<:�}g��gg���'�;}U�@�,�[Y;j���u�����VP%��7U�RG�Q���O�uĈ��[��O�`K��[>Re�n'�W���$��7���:=��E_��@�<|}�&w�})�s����/�Z���϶#��J�����[|;��#硜'BΘ�*
0E�-)̭��ti���o��o�1�IB���h��yAp_t�g�C���*];7�=s�x���ecӚ��o��[W�$��%�����g)W��$`Vm�C_nۏ�n>�]�g;�t
�1��gOlԻ���K)�0^�^�p�Щ�[hjg ��=�F��S�f��_+Vo��1U�3sZ���8E�^���4�;�<��D`�W�\B�A�T���b\�*�x�l�Q�{��nj[�~�N���m�s^�^�l�����t��{8����j8�����6�~�x���q� �~����"���Ӹo�M���<dנ�8��yછve�ʈγĕ��p-�X[���!�����^^�b�`��\�}������Z��٤�`˚��|�qw<�&��\�F���b(�Ye�ig9��q��̢��+A���U�R/i9I��-�˝I�n�U��Cq�d�fC��ݐh�2f����5l܌*2�َ���8޹�Ό��;�{}�xC�֌��$����(쫩�k-��˨g�֭h�.�os��v|�{��1���������9Nŗw�+r��ԓ�`�p�,*��V��b92�؇��PGC�SS�_!�^���~�S�[g�f�<>������`��Ya�;{�}��K��k��0,V�&n�j8$�=�'V=�XY���m�Y�_��nn {�N@ݖ�-����]�V� wP��I�Fu�ˬ�<_{k�=�݅�7����=���GOw�����N9¼�G��V���9Ǟ��rd���%���5š�v���KS=��s�Q3�0C�i�xe��!�v����o�y<q	v�({�G���o���͐] ��FU+����ս�zvI��~3���~��t�hӼ2�I�ٔ�p^ـ��b�V�vk����<�׼B��ͶKrt����jc�g���=N�����
f;;���睞G$=u��=ټ���?f��(���6�zw�za�J#�LP�o�[�����L΢��s��5Qw	<W�
}8���u[������Թ =��fnh��n�r��%���ov����[�\e�p-��C6w{÷�̮%9��Њ��x/B��9NE���o����Bf�A�El�����"�P�I}%�B��� =�j��H�Ud���M�]�vY�	����MY�7r��Ａ�Ci+r-�1ލ�2�ЃӁ�����o�ɜ����zx��n�34ǅZ�<m��F����n�2M��sT~����ynF6i�^V���;�j�p����ۗ�����/�
³��0 �X3S���sM�[�zk���|�xH��,9�u${ڢ�-�JvD�	I�J
/�G���s�"�j�yP"4�\�x�3,��7g��N��+�L��^����tIil���46�o)vm���99x�T�1�t[aߴ��]�[vT�W%:r���"[�ݨ8�X�;���3NQJ�~^�%g���^5��0��>/��z�B;U�waP{|��V�^���:�dQ�g3��ʳ�7�����o�G������۳��˞柕��gt:֊iM���g��/k#8a��0B�~���{d�F���3����'��8��6�o�:l���;�3ꗦ��ާ�{�;�N)��I�nW��:|�K�{��D�w��a���o��<����el�{�ޙn��]s�[@GW��^ޫ�zaf.�/���A��$B�5�3�3`�w���H�8x�OJ�����=���� �<wݻ�Xz@ɳ��;C�0]K:�o;�ZQVN����m��qz;��<�߷��m����W7��T��6�������Ho�����6W���R��᷻��z�{��yY���v�|m��=����u?��3Z���k��;�H�TU,K)h�o<�y���^���qڼ%�����C�(�g��4�G鱑� �}��^u�t<��$ ���֑�U�j�듃s8Y�T,�������2)1/]�pfS�� b���jSZ���+�C�[������;t pWA���އm�u�㞉�vû�z�@mtNy�z���1�Xx6����uͳ�ŻY��hl �A�B��]2l�vpvZ�\r�
�@�u�7O5���;��;Z���Y��َcA�yv���ѣ�ڐNr����gVݵ�c����%�7�p�q�v-�7PK�n;V��)�e��g�x��h����f�sqsgy�:��3��v���rvk���<1���h8|�Ɏ��l��6wV�OFH��O�E�7��j�8�ɔ�:�=�J����v+�����ː帲i���٬�7dݮ����`wC���vnwl�k<�L�c�5�n���:��7V���s��c�qW:z��&ώgc)�9a.^�\ȯ�Н�X�X�=;���=���1Bv��9]�s��Fq��������[9��,/k�����N�����n$7c�n��d�}8u=]rF8�Im�.+�W#�y�s\f-�%��Xn�[��c��n��R��x�?�㾴�J6��� YdC��q�˄�U�4^q�s����6Ϥ�bEVKm20s�f��Q{�qh�	�:���yF;���9e�
�w93��,��_n���8g��rq1� 3_a� �F�`a1S�m�����	�N�į�t�E���$ar�!%l ��	�[r P�v�d-#԰�|3u���Ul��Apo�z�D]��_��]�����V�ߨ��S<P��WY�(p#�'$=���F�K�3�f���`��r�h��5�&E@��ϛ7�,jXQ��E�)�7/[���ww4�7j&�n��|��e�͐�B�noZ�APdDtj)t�*T���lX%8��5�"d��*p&�)�L���^?/)�\��3yV���d��Z��U�T�b���D�q�vWٚ�T��j�|�yY�0�z֌乎�'Qmr[n���d�{'Ym�/m<�y�1Ӷ"�6�Oj��l�h������=�^��&9��K�=��tk�j��g�۳�Z���]F��ݙ�����MV˰<ӧ����2��M���e�U�շb���¡�϶�_�����ߊJ��������}�	���j�f[vLe`�ǅYm$T�o0�/���(�k���\��Ģ�ޢ݀�0���i5�+�� n��I�`��6F��l+�@۲���БuN�z�4}o��梭�W��}��U�����sݳ8�<��hm&����ݞ$�b~���I̍��B�O*��ɺ��� 0<`��lޗ��I���0
���k.éOt���w�rp�y:���9�z� 4�J��)pi��;R���3d�jW���}�|0H�YH0er�䮻45�M��ܳ4�YV�߷�y\U��o@��Ԣ�b�B��(�7�@�¢zۊŃ��+17��)J�b�;~�����wR�f��#dD�P�p*��a l�v�򁲢�Q����j�uj�DB��;05u��Uf̔��
��&�I����I��l�kV�gweR��3� �l��AtU��Ò�{qm�*!�)��Z=z���}Mŏ{U��b�L�1h��瞗nh%��L�ťM��to5t�u��]m�ë\Ai)q�W{��\��AlU� ;잂Yd�L�rQuO����*:��Ym$T���ad^5ԓzI�t�#�3� ��t�{[�[$�]�oVg.�P#��ΰ����~���~=�JЋ7��"��DG�wTe�֓)�(��KG�̃϶\��c:��r�I�U-#�TZ����`ն��؊LR�ؔ]�U��%Uѓ��6f+���x�E��8 �;q)l6���6s�{���61&H(7:=�x힣~:�^AÍ�.!��]�N[�bkQ��J{hv�譮�]�vY���*���ltENo{|�L��z8t��6>\�WH'mf:�V=:��v���9�s�O	��g]���B'E]�a�+dݬݗ���!�<����C����T�|��u=��=묾�Wn(�Y��uv$ר��[]u�|wۛ���SL�ɸ�8�X��Ƕ۷�m���2e1Y�oc���9��D�V=�EU7Y���^��C��I&/o|<�/Yڥ`Fnb��&QS�I�������]v�0��R8 �Wg#��� /�V���$�(DLWcq��$g|j�Ėv�զ�4�$�::�+��F�)iWb�v^�������7�A{R��"Z�$vkά�vږ�O)��&�M,Jx�Jw��M�̗�c&��]��g]�@�6��|��&	�:�����]=����癇V���R�
���������A8�2����j2�԰ w��="��EL^���3������o���,%� \B�\h��[�k`nR��)��NE�jQvC���"���2D���f��xUѕ�������h����s�d�˷}���]�b*a؎9;�&�pv^����]���$�("��G�=�x�҉��J2��iΏ۲�5�+<g�fM��ԓA�bz7����(��Y�A��)�IQ�QH�+�)�U�u����������f����,<��k��aE�1ڻ�3wm�j1ZVx�ц���)'1z���r�{�q��F�(\e$���b�}��o���ECW1|{T���\�R�:�N扊�.���M�5kξ���8���� ЙL�"2oMQ��2SP�R�ҍ��cq�m�����ԑ�PU�B80n��:����%h&�����u�Y���ux�EnƧ���;F��&n5�*S��&��!L("z7�ʶ� {Z��ol��ZEI�x��rۉ� 4�J�Q�5�e"�;P�=��V�ۂ��b�Y|��,��w�6M���K��[�$P���WtN�l2�tUeG��u��5ګ����� �*"�U\�֡<�g�m$^�U�Y�v���9��m�;sO��ͻcj��\��9��Н��ݮ�GbN֋F�:���q����oc�ݺ�˹mڨx���+�q%��c~��4(Y�^�r�����?]`��B.�끇��Хg]Е���WjԨ����y\U��o��Ԣ�v$�a\�ՠo
��n'��9PYmە٭�b�{1��Fgb��)"�N{چwS���[Y�{�&b�t���)�v�|=�8�ێ� ����ν:�1F���ղ�F�_3Qb۪�/f�-<\خ�沭��]�3ي��YmG��N3I2�rLNM��3Wl�����n�Wj������H�Wy�Q2͙Gb��n�;���=����a2���h6�4ƛM��z3��^u����.9�"��:���ӴK��I��G��Դ枳���C6.�.	������p���*�X�Z�߅����	�W,l��Fg�:ۅ���`e�K�(�J:�}�x�q�X�E8EDLWc�zM���z�%[�I�$!�)��n�����Y"��X��܆���z�lep��8�e���'�"��uMoP��:cG;M�r#�b�}Ǹ4�w�~=�Rj��3��] �=���o���sR.����_LWpD�Zr���J��+���k��;����>��`d��#�@�Y�{���ٵ��n$�����X��ݧ8�7@x���}��Wq�B�� h9@<���=��c�]�����G���Vg����j7����B>͡u�S��]�	��yzX�����������~z��[���j#D�Q�����3�W�߻�����jrA:�:v�q(���Q�J����3����A��7A�Jͬ�:�NƺY(VPGd�0# M���){{�U��|�߰<�ʑ<��s�ڗ���15m�_��[�^>��� H�&�w%�Z��`	x�?��w+#Kp��r6a�m�3E�K�,<z�����τ;�~����~���I�(z[�ݸsR���1o5s�Dad�z�w;u���x��nhR��Zw�Np�/�A���YD;�xBKXp?���E���>�{.�����+&	 �=Aؔ���x�s~D��?z��l �qs8��e?U��Y�L��9.�-�����Ü��Y>�bѡ��Ѻ.��-��t�� 4�����oF�T'| �[�G<� �p�	n���#p����я���@`�;��W��(����YMH-�O H�`��U%q�4�T����#
��4`��Q{m�@ش����8����5�"�������mSI��x렕��_��{e�v/���ļ#p^��pӀJfR{t�������II)0�؛llg-��u����Ktc�]���v%Z[�o�_fS��\$��q��DI7����_^u/�g�l�r麍�x+�1���]\nGG3���I�x�#���뷬�N�����A��="�����xw����j~��o�,�Uk�e��55�EA�=!$^=���Yyxϝʒꤘ� �{���J>�mh��W�����aK��ܻ��P�������;��c��	�G�y�瞐P���dD��+�1��A[Ø��������rG���I.�&~}�s#�ǵ�����h�22�S�HF�*�hb�l�:��X��e���w}�Tw�������n/�t���T$1�O$y$c�ſr��9�F�K.����Փ�p�d�� �B�5���d�
{����J��n���<����q��A��,���܂���{Vm/�(�J��*��U�![�X����
Ȫ�ު���9G9s�og;�왍�t��N�谦Q#�N�4;	[%�]pr�j����gu.�'\�w>�k�Z���d��;�� z�۵��s������ֶ��4any�f\xlv:Ĩ���jޅ�	��{n�ܢw�{nݽ�{vd��e%K�\�����~q���O��;+.Yh8����I,�-�t��ێ*/�w��2���/u&JjJW֗w��ݕf7zV�?/���!8E7��zG���.�{;�u�1;�����m���;�c�m�֑�
���>{����f�����1��M7�¯ZG�iWK:�H�מ�Ѻv���TW��3r<�Hfͷ�ҳ��_{���g�5��C�!�n��Q[1��(��;�˕�����`�������4�[����.�Ay������#� m�r(��$���23`xF��fL�oy����k��K�(oj��;�6#�޿���=���j
I��x����r���s3� y���,�mۥ[�6����Q�kqZ����5}��E%�Q�وRW[�F
W@�Oaa+����[hns�n"�����|=��Y��K3�����y�s�� ��9�S�]��q��b@jl�i�lğ�}*kw�H�t|+f#��7TEVnD|��T�\�nv1�7�X��&�M�9��4���bF
��\q�	�m�^ϻ+��1��N\��	2��<$��V�ə'��{����ji{��h��?sl�����6��o9�1�- O�?Gl�Os���*�s�ٌk�V�r��K�� �m���e{��5���ڔ>W��h��Fr�� ;�u�UI:��������L�m�)R���s�x{�}�N3�C�ݶ!���L���� 3�0�Ƭ�*����Qs�1)�O�v�<���J���o��Ь�~I���W<G��/�� ����I1��� �Ǜ1�=�wVKm޳\��0��>��_l>�>a-w��J�J�%��)Eh�T"a ա(�5/�O8�:1-�i����[�����|$^��{���?~?!A|vl���,{�����I�a3u[�T{G�������h�$��3'3&pxo���oOQf4�K���L6�%u��������<s�M�l｠ <������-�)'&�2�xp���kL�6��a؉����Y���ر������OI�M�� �n��@�TU��w���k*Q1K,dl��j�n^֚ͷ6S�yls���ƺ�(�qR#��T.q��nz�p�x7f�Ft�n�Av�t㇄���=�+�T:���zHz��k�b�nk���k��YP���wd�#"a�H��P����'\����s���W���{tmR�~����nL�JY ��>�'8�{��_<?�]�<���LKE�2�����{� M�0������y�����;�J,���?{�{U�^� ����׶䕊�j�rB�%<qHION{W������ԁ��b����rQP���S�]ׅ�$�*��F�]*w�+���Pǘ@���*m�F����)`;	��1��(��W'�f��d�.��  �F4�+�`�d2�.�F����ru�b
���������l���}}gdoT�2b�{��̜���8�4���llLl�Bi0MM���6�$�}]�/ܒ��<�D�cw����[���3R����T���L�z��2[���K�c�Z����U�Uh ޚ����4�FQ�g� �{&$�s�S_��/��\(i�W;j�m��k��(^#� �2�"�Q���̛�3~A��ܒ�}�X�ķT�^����^q�O��?UΏh ]��]�̔�H�6c⑻o������Rm=�W�է$��22��V�]%����n�yu�K�������νy�{�##6��#Q�͋bLl��",b�d,��~m�_~}��G�ܩcB��))?���S;�3&�8}�{���T�٧��6��qG{�@ y��>-���=�t�$"��s�J�ώ:�6]�WYG���3�i)m74�|e�>Kg���x
�uGq}�2�%�J���������l̛��{���U�tŴl�&l��I�R��Ic>��w<�5O����N�����}w'~N�)CT���#�����{���2GR���fA�w>8hS��;����5�lh�z̑Jlh@$Ţ(K&�b�L�F�h�&��Rl���{�����M4�A�~9ҧ� Ψ���~���������@~q��"�۞L�g-�z�����ћB( ��Kfv���ya{I+��:T���Ȳ�nI�[�������2w�I�V�#����݃�p��F�Y��A����˷��m�;$�SH��ƣ��y�3��v�����e#7��B�1���G�Y�/�[�{E�hǜ���gʭ��T�+����:e��g"�<����}줁�<"�;}{����w(AN�g1����?E������i�dc�W-�#/6 ��l��پI1�*-�5��6=���k�V�"�r��k/�ë4*V�LР���x[��	���xvĥlkk,GyU�0W�2hc�f�4�o��w=3�`����}�J|	ñl����0w��1�n�B:X>��̈́;Ȃ&`d
�����ؙ9��lrn��h9_��q�(�w���vHtz*����IJ�q��,�_�7�Fu���~ݥ�'��2;�@��X�����uf��;*�g�{�����!��f��=�"k�ee]�1K����C
f����Ş��_x��mt�u�K�T>&{����ofr(���*�&�Yv*��E�	۶�> e�ˣ�QO�J3ٿR�Ŋwf��{Z�IGN��n�/�MU���p�gWv7I�u�ηgT(k��=�sJGf���M��h$j$MB$�;Bc�u�b��c��n�g�0d��"��\�B��۞F�oh4˛Gٍ��l�����@�0��mr���C�N�p]��F)6���ss��A��Z���.w�<InL��L�T���.�܈g� tlcR÷go[r��n#VB;m���:�۞ܛ�}��,��`�l���^y�[k��<s���ɼv�V�C����{V8��Wr�tc�M�/>�v��1j.�cF��'�۴h��G^:T�ц�v�0\&^�,lU��t�s�xiU��Oχ�Kɚ6�ٲk�\Vn���J�)�5F�Ng���Ƶ=�@��F ��=u�f��!�����U -6���Y:L]�5�[��=]��u�N�4�:3�Y��slv׫�3�N fG;Ż;"ʃ���6�ގ��rs��<&끮j�z�[qk��2`g��]�Y�ؒ����8n=��n�l��7ku�^V��r�r�%�zQ�r�a��� ���a%�v;
(I~�c�~M���#Sң��4nƝw晣-RLu�oyy��'r	wx�x�m嚼��t�ws�;X;5�M�_,>�y�g���2�d�M^�$�4}������1�7(]MBoZ�[Uxk*a�e�֗3{�r~KwO�׵Su1��p�H$�VN��/L�N8�g�.���L � *��M�d�-���g��H�m�I{1�C2~�6G��Vx3�~�.v-ҋ��E���qx�ۗ���r|�������%怛�ɫsj޸7NİɡL�gEgAG�;�̝)T��3�n��)�����C4xQ��/?E�nm' ����E��m��?B��E'+��e��n���,���4��W�巙y�a�	`�F �e3L�m���F�xT��<��nr�D�]��93#&�gyڳ�qk���+B��U���
W���tC��: `��q�7g��Vq�x8'[n��nlA&/n�$�m��c����nM���Mr<;�� �q���s���=x�玵ǲ�6�&��x���v�v�����{�攄LBP�B(�L������P4��Ӯ��/Hi�7:�GZ9���Р
)W�	f��Ieޮ�܌��#���=�x7������(5
x��?x{�Z���)��{8ƍ�����F%�H���Ҧ�w�<<��~ݙ���֊E�j+�� ��5�3$��- h��jG����))'�m��x}�xn���}FG�l�1�.pj��h�
�粴
�v�K��{�%��Y���#f����_� 
n��qc�$�,��|����]Y�9�rV�S���AMo&���N�ڻgW]Ѯ���I�(�h�1`�R�ɣ2�"S� �Rl�l�R_"��<�����h��*�-���p۷2w��5h�h��fV��G�<�y-|o%M���|��}ɥ�m�To�32~���j+:�3����ָ���P�J��Ln燐&j5���߻ܪ�:��ú$�����������1�or=p�W%��9o��< �^y����s�p8�bI���v�U�F��kZ���[�E/��� ���\y��L6�.:�I�J��^���k�i�Dx���+��5��cj0cmck�xԚr����i�F]�S9�8��'�N땾b�T����==�l��Q�P[�eB���5�l���s'�vwY�m�6a6;�I$V�*(Ъ)i\%@��1����4pSe��^o�Y3����� z���X8w[�%LW��xw���ZLq��ʚ���{}�y�{��(5
����2l�>B�1�u�I+w�]�F%�������WY�d����.W��ݗW�ɵ�g`��g������s;�2�n��^���QX�(���� ��;��g>�E�j(Ɣ����:�sU�u��x��~8��BR��v�h�rq�iRv��8�{��)mA*���ٻ��7˼;�z�ґ���I4�ITO�����)NmS����{�%�y���������[�<#�_eܓ��5K�i��-�U��s�'��~�����ޚ����QI�(��3'���>�~9����2Rr˫������:t�X�W91u�;���)Lr����o#C1f���.{���%ŘY��I\�U+UM���I�P�{g�l�u��q�q���P:�t�࣎�Iu��=mh�t�=�s��m�5i�����չL�hv��a;3��-�7Q�9���p�k���C��5�0͌Ew�;<w�]Ȕ��N�r�P�
��6B@@�w�&�FG��}�%�̙8~�%��I����}�zo��3�>�Ա�,cZ7���B����~���g|�����a�6��|t�S���âIc�֥ksX����RI){�]o۰�2�"��a��{� 5�n<��$� ��.>d\�(�cTVX��pP�ln��t�+�0�0��r�16��;��1E[S��{��x�yG�o���;uu�@���ڟ3�֯�q�A=��pX��Y����S�ޮ��s�����מ���7bK60Scccci�� �ֽ�J�d��\�}� 
����CL�Q�sq���K��ڟ��I��l"�Q��{�����rw�ᘲ��o� u�]��ܔAbO�6WW� �����7��̩�X]�u��͡Q9J
����5	-����p���-��N>G��oCd�<=�yK�*Lg��M�IRO����Ownd�'ŕ��=/�ϖ4�e5D�0���J5fG�U�M�=œf�7[��j�]�8Q�=I��sIŗ�i��s�]�s�y�>*4��Tl����61� ��nW�$�^gn�T�
I���G���3R?So<0�K-n/�&SE�n�}���� ;����3&�6yc{�<EHHV��Tդ�[k�vVYA���a̎d��Bnϻ�̓��?��;�V=m��܉�S�|٪?n���x]��8`Ɣ��S8ot��f�/��J�Ǔ'��?����fd����Cu����;y3$�0�&�g�g�Ә{�dп�5�7̽H���Y��7�>���IԈ�= 0RD�*�����μ����e8S'��~���ٻ;��N� |����b9+��J�:�Ylr6�"j}�f�w(�-��n��5�_{Ç���Ę���D������da?U��txo�+�q����&�����K@���)����s�j!����~ު��*>7e�4|�N����)�1
����2~�@���,rH�53&�gEl|��'"��~��"�9�(:4Q:mϲ�)���ɞ[4(��ʹ���=���D�i�̗�F�	���A��c��"���k��K1Yi8��P�B�Nm=�SsU;�j҅�B��خ�v.�+�w����f<�lў�m�۴�2;����7W/|X���K�;��㳷l�ĸ�m��:|,bX�ZV|���őW#��}����,��^>S��̞?w�$��k�c�~e]L���:n�=��G�>V�J�K�c3�7���C�?M|���EU�����C<{�O�m�
;��f�?�L��I97�d�0ve�&d�F�V���}ۖ�u.z���qe�kuE�+L��R�/>~9�'��~I|�v���9���$"�r���U��;8��C�q(�ꞷ��^�d���]9�r��N���|��ɰ��m��m�6G���ьkN�)���{D����%8m����LɽN>���Pٔ~���Z��(�d6b{�#À���=��~��w�۷rs����a�n���#����wd�1g������/�E�	�j�����'7��ҕ�E���k�>&�M��ͳws2o��*�=��*��EVZ\�{c¼�d�ʟ���`o���6s�mܝ��I
�o�:��2�]N~B�v.ܰ��������|�=wU�yf���y�5c5Q)��z91�.�dꉕ�V���,�b���|r x�/v����W�\��Fȸ	^�P��B�Vq��@���u�J�j/2A���q�XN�J��Ss��e�hc��q/�n�M�"Ϭ(���c-Q7��h��@��U�����q�5~v(����Nfݑ�T6�\5�Ŕ�U����̶�Q�W,~�P>��M�z�_,c�"�{��U����/��	���ھ����&�N(<���T�����������m^�����s�*a����K�cf^B�B��8f�;�&d�z�jb��`،���V��}�r�bt��e���ws�;#��IX�4�1�70,���娕'�b�llIcM8b���Ƀ�"2��ü������D��่������Ӱj*.Mx\C̵m���M����.ST�Ł���\@�����l��M��e�Tz�9z�̈"O�h��Q{���E����4Z�h���U4Dy@�8��M;��u�u%(�*��]��Pr�DyΧma�Ҋ��ԃzR��>�b"�@��T�9e�s��V~ �ݛ��r��������B�JZǼ'y����o�R�lCh���+�1�t}�r�0͘s&r�'��6���A�ry=E���x^����sFo�4O������sՖ������ʽ�]v���l�Eټ+,9�j���D�b*w|���jh�T�`�[�)�"����L�e�T��!Q�%�Ϟh2qL ��w<�u��ך��3F�{x�&�M����d�F~�b�78M*U�{�GuU����gG�����Y�n!��a̵�੓���LI��ʟ��w�ّ�����哧�]5�㞂�Y%g�fe��q�,���LɽN����/�ə$��H2~;�_ &�L�k[/�+|.���nͫ��l�\�m���<weMG�>R�I'��g3&dާêk�����u^+����hQцB�a<n�r�/�[u}C2WN�]Qm�i�1���c��n����WRT(��yG����m^BE-��w��/��n.w\��#�lk7#��J+e+9L�HAKi��Q�v��u< ��Z0��?�L���U�Z �D��6{홓|��U�����e4��z���c����R����Ƀ'	�U�� l��w'~N����uFU�Z`�P41'�*{޲�k�e�왒K��]�Q��Fټ̝ˍ�6�n�aɜ*и����t�S����
�_tL��kk�6D *j:X� ��WX�{:-��9K6ାy5Ѻ�\Y��OZH��ך���u����uH����|��۫m���z�y��7��Þc���g��\�9��k"�󽷻sm&�xm6�efb����h�ڹ��wJ����Sv�s�Ɇ����753$�<kNd��#���p��7����2w��)-wّa�Ci����a7r��x^D�;��OP��6�s��Y�a�����fs�%��3��bna4�U�D��2w�fM��.o�ZRArBYH�r��ca-tqE%(; +d��=��2N#���N�d����$!�*�۬��_���䐥�`�ۖ0�c�	�0EF�mJӝv�+R���=�!��6��L�3�f���9&/z�s�e[��0Cb$�_��}[�dπ��U3��̞?b��p�5x5��3ٳ2I�8 ��[��1�S)"������}���s��#��N�ko窾n"',�u���NnB��wC.39��(�YE]���6n�OYz ��[f��IBp�)9?�<�(ґ��fI�s������e����Wql����!�u���<�npWmv�G+n�����+��i�Q6��Y�]��VJȿG9=�F�"���` � �ovVϻPV�/u�I�*���?>��uG�w*wñL�w�48@��}�3��S��c
E�	�%�g�j��RFV���p���V�0��9,�#�����,�Oc��L�왓{��L5�Q�+�
<��6N��m�xM(�[P�#$�6�������f4�z��A?4��K��b�%�BD���BV�p�vf,��s�n�Wpqm�'Tb:sU
�۾g/]��6�i�m��1��k}�d�kk�;3|�=��93�$ݎ��yk~�MIa��-*aX�U�t��WMfkԿ���e&�w�{�Y�sS����m��W��)j0�w�.j����z�8��1��}�̟����#ԣ5K�J#j*�`��"L�=�K�1ԕ�Ǻ��թ2�I=�p�����[n�OD��\{o(�WTj4�H�3c0�	ø־YR�=�����s��L��Wc�y�*�k\�Y:��\�������lV�]u8:6�v�3P��9<3�� 듩���ǰv�㛲�$3؃!��fwL��ڎ��g�$����BZ�Z6��;뮮���Q0�2&�t���Hf����3z�tv<(��EJ���YJK^�9k���z��=�}c�RSl5b>����vg ��Y�T���e�I��N����W2��a�g�e0�.s�¢�(ަ��7�+�g�e4���U�<s�{��9㏩-h�ۃu�K!%�ѺLGh5oEr��
wX2�[�����ᘫ]�w���'Jb3ڳw]���zu�3c���/e{��]�����>={�1̯L�P/V���Ѵ�1�(���ۏ�:�=O|$�臨��6'�}*�.��G}����2,��4xWt�ʼʙ9���7�Y��4���I�'��x{c��ۻ�@��u%��{J;H�pŃ��gN��U�,1��Ւ��۴dz�	�K͜��٧�Tt�p��Kv[7�3'��< 5V���2�6�T�kl�F؇����g��)��)�p0�86b2�N;/n^7�߮��z������^z����D�1,�I��xI��|޺k9��Iۮ^Q�BI�U��<��?��R��
�e�V^ ��p�1'�ٙ��^��{[fz�d�X�N��`Kk%��d�2�
����8�6�KH
�6�}[3M�y��k{&f���e�H���ޟ���I�N����Ҿ���)��TO c�ʚ���̓��4��)�,$��f��b�6f�g�x���JT�+���<toWf�M�y��&��T�]w뾺����QL1l[�֘Fo�ęL"��Z��:�fd�d�f�Fw	sw)�x��Q�1Ul�e.z��w^9��rL�+SL�6ɴb7���j5�݃�����}���Ky8f/fi�q/�'
[f$��35��yv̳]�2k�C��n���GyK;y3$�0��.̪�Ǆl \&�����̪��t9�1x�ʿ/�2/5����L:������NO�tlݻ%'�I���;ڣ�H�}헎��X��
���܆�>��&��Қ�}�7�8�t,E�i^ë#g\�n4�`��6��Ɏ��DU��M1����q��.�d���}U��GBp�.ZD��3��=��W��n����{���o.����lI���Z��5��tT�A�j��f�ap��m(h��q�֘@�j��T+�'a��Z����3�X��c\EJN[#U�̉&wg�ڷ�Q��t��x�r��t�ÏӺY�����C�fo�Ws�E�n������1<���|�_�8���|l}���rt,��yW]˞�yx^��>LC�I�dw�f�)I���{aE~�oץuk�.r�"
Nb� �w�"1�x�6��7Lءί5��ES�Q�N�3c=N�ʿK<lC��N{��d%�ƈQ�<�7�މ�ξ=�-��u'Ǚ����ry栙�q`�����t�Չ�\��%���2�WL��y�m���ģg83n��e��s����;7��8�୑e���(<Q�|�z,�W��ױm͸�ݸ93�<�����q���z6��[<��9�܉�cr�!���軱ci��9��ӷ��6y�FM���P�\'�Gmҽ��B@�Z��J�z��v�l�C"�Vm��ع�\���kk{ !�^���v��� <����k�	y�7<����=�'��x"<��l���m۷D��Z���tSa �XL�=��K��.nҗC�OX���Wn��'g�H���x�����g\�>{V3v�P�x�\�\g�^�[�/d3p�v֋v�n)�Xc�.���Y���Ή0���:������]��u�(w\h�r�w#��{��L�N������.ȴ�B»l��;)mʜ\ݺ:ۮ���fs�\ܢgr6�H�����۳'(C�1��v�����u�Fp�#��z�a���6nv���q��kF|��$��.�RX��۞lvjj/n�ԛ�v�
j}��-�[dM�p��=SНzc:n�j ����fq#I�t��G�D߅��m�x�q�ܸ��=��q2�m���x��oH����hh���o����{{�꛳�|]=Y���|9y��ͱ��o6�*Y���J.�d�4 -����<�܋h�3q���(�%���G�e��O_��&�4�ǽ���T��b�q]����EaTf��E��ҽ��`�M\����By������oy��Ε��3��Y�s9F:I�/rm�5nۜU5)䴁���j�N�%�Z{wt�2�mb���H(��g�r.Iy���R�.���AQ��l���x��X���v��ӑ�Q�97,�2#�d����g���v��>��.qto=��Ϗ6�8�v�y�pN�^�Bz�Zͷ(]�F�Za��!1�#��X·�u��$�������=���*5\qcRA�~y�s7m�;��"��1��u��tu�@M�!���������,��I���1�37�c	%֒m&�m�m6!�ҬS��Jb��\˥<�f6�m��f�6Z3����쩟��`ѼL2�6�R�y}�U$�0��s3��̣��jq	C0aU홎��3|�=��9�Il]�X+A8���ȸ��Q�>[-��T3��"LQ�陨���}�&UvL�Ӽ�&[	#QF3SЎl��l^�+7�iŵu�oV��W����{wn� xy�GM6��)5�oW����w:�EoA,�	BR�jSvݏy��/��ٌ��e�Ǒ�9�35��-ٖmw3,�Ki��ѝXVo�$����;8�����&�b(E���(H�M��H&�R��o;��Y�m���K58y���i6��V�JX�#��3Q��<θ� �����2o�w�Wu����� �ڭQ�dV)���Qz�(Y#Vм�t���Qs��^y��%��Y6��c�MS3m�ԉ&�Kg�\ }�T�sh��������M�D1ɦ���cy�~��&d���=�LΏ\
�( �G.��i�0[IY���.T�sl���T��I���=�i4��B�'�{�-^d��kh�7���Şp vg;F-lF�^�g2r�gf_�0�a��:��̳��5�35郢����[��3szY�9��������]���3�Wc�/�d~����	QhL�M�m��3y��NϹDK2r��=�^����2g^�={��'��1J9mV�-��+h��{g�=R��%���w�̟��ċ��m�kY/`��"LI��g��5ze���3�9�*����2�I�1��9W3��a��s���U�Tx ��e�̙�|�'��sT�v;i�["���a ̧W	��/�i>LB�9�F5c��Uv;U���t����ú���9�zc�q���Qxl\+U�7R�L��ۈ$4��ح����s۞�n����`ĘVj��:�r�i�Fu@�uWY�DG[;ׇqe��n{<��(\�wWR�a�ֵUTk��\76�x�M��(q�8�0�us���x��TIH����v��yӷ.�\�ݹs�\̀�n�ֹ[0��a$����&/g�'���F��~I��4�:�K|Y���fM�'�s��iښ�۵2N�� �-��JUN�$JL�}���Z�3i��Us,�N"�ى1��燽e�{g�\̜���҈
fL2S{<��^��6;	��=:�,��l�6��{���.~_/�%�'�oNM��6���� ���Y��+^��������r���eMu�̼V�w:����>���I40���͡�m6�������{�x����Xi}��
�'�auwS��f%Sy��9�x氮3.]ZO��£Mq���i)��p��m�Xh��ެ]�g���v`׫\Z�/9��R���%�-WW��7�J߷}����6��	C0aLm��� �;��ás�܃6&b���M���b)�z��V-����N����@���������!C�gݽ ��t2�-}��Z�QEBA���;5�c7o5�ήT�����]���=y3j�~_fUN�(�	G��x]ʙW��1��7���$n������v:�2��= ]N�q�Am����*#.ۚ[�l��پ�e�a�ާ�xʌ���ə:V�x�Ul��k:�@��w	f�y	�Q��&�
iڗ��]�/t����z���o���>�8���m}�m��˱R�5Z�11y�F6k�S*��Q;]x7b�*<�m�cEF4�BHh�M�󞯿���ߎP�+�:�x�?w�l�Q��6~����|ϝ�V������5P�U`;��Q�*����s�p	��Um�Y���CuQ���%m�L�*��U/wCQA8fd�6��x �z��*;Sg�݀i��u\<��9�34��̙qy�L�j/m��#�������B0*
���5��xdo`�/!T��re����#3���8��qh'���{�.�r9٢��J)*�֚!!W��z6��!/�]g�fy�SXn+sF�M=s768�n�өǢ��k�q��t�0��z��!Ш����N�<��{Ȝ����)���Vڭ]]���A�7/M�W+�i(0�h���F�N5��c�Pl$ʊŞy���fpi�r*�LЪ(�Ej�dT��;���-{ݯ���}�N4?ja��e%/ٵ\<)qp�ٓ3IX�kb��%��T{[f�8��Q�)g�&d��f(� .I��{�u̳�Nj���j(�jl���UT�u�=���<K���l�V*�B���<�ݨ\$��\q�"�!�sl�6�j�&Ln&�Ƀ͆�*��Fqˉ���weӳ�u��^�I���Է�_����]y���ـQ�Q�Pb�$EE�Mc��B�W}������H���	U��4�L"\���d�M��l�۹'��fi��i2�55�m����}9P���=���I�[jY��fN���=��Uz�:�����!�hfs8���F;CA�l�wg5�j�f:�x	�ד2s4�
��I���{�V�=����	�^�Ɩ�jM�M����1`�SG^���0�_�S_�{�����wC�:�-ձ: -J�VC��/�4]݋P�� �~6��N�9�9���w�g�>��(;V�ٍ��ݷ�ޞXZ!�֨#��ŃǞ9�wx�q�<3��M��otܙރ{����7���8��>�����wi�z��N�7����f�e^[��9[�Ϻv�8-�cDMG�_�����[���գ�q�0�θ:9�owY�s�Ǹ{q��L��co�k��:-��o۶���e=���T��2��������}��}w	8�8� u��@���0o�Mn ��n���9]ނy�|����}��lz��~O;���~���u7�c��.��qdC6��#��.�&{>�.
���w��0��a��z?o?l��V�qɌT�s���=������gSj6<��ڒ��	�N'�p�D%{;�葮�"�.oM�4$��.���:��@!�;�m�2l���-7O�������ﮆ����C<�ol��0�7=귆r�`�<n�l.�{����K֦�n�Rr�C�B�c�b�]���/��}�ڽ1��a�5�ǻE�E7ݗno�l�$.\���h�QZڧa�ys���OjCF��p��23(���w\�-�b���M`�u��OQÓ�t���V���2�[,(dj�Q�K^�I�s��,� �Ey���t�sI}�mڔ풠g���zv��E�RR ���'P)0lSYHF�1|���ˬ����LF�Q��&(�
�ݭF�۪4�hCIA8�{��g-�~�����r���v`��'1� �#��3�U>f��vQ��U)����+�u�j�[g�Zx�+Ci3�jQ7e�Z���
Dq�X�"�iK�px��i)�~�}	�)��JY�ٙ8P��5ٕ3d�V؄�0�<<w�^����l���Җ�躚]y�5]Z�\N�&�\s������n���1n���}�p�k���Wގ�$���ě�#	b(�ɉK�X����{���}]��BF{uw�Z4G3#�n�_��LD[N3q�Ԃv� �;��
A-/���緊��_C������ v�x��]V�)�� �2��i��3\��a�4]p��q,�#4{����uxZh�-���E25l��qe�g zh�(�#-��-a����b�.�u�a�|�;K���\0�-���Z2�a"`�e��?J�)s�����nQ�������FYmwx�a�jؽ>���'7��_m
���ݺ��4w(q"��	��]���4pT�&T)�쫘ݛ�f�n�H�kn�8*�(�`�l��cl���X��޹:k�9��[]v&� �l9��U����zݎ{�^n��[n��Ws�4�^;E'<s;��n�7-�U�gy�z�t��>I�Q�,Q��1A��H�`���?>|��o[zY4�⹩W5-U��±�����y�/
��w1e�,�����V�5^�!�=3-i�r��h�kX��rUۢ�Ѧ[^�s��3MF{���5���rᆰ�l�����$֙���-ӣWu�S2ղ��E�a��jQ��0��)a�2��w���-[4��z��[�ZfZג)��Z�E���b�FYm_�Z)��I���Y�x�õV\oZ
g.��S�Zj�ovF��=5�R�0�.�ˆ�E���>���	��q[c ���
��0�"j8����X���U��*�L�[+z�Yf�F��Xh�ܥ#-�^�~��[��afZ=�Q��A�3�v��ү�'rk���әSpL��������?O|  � ��2YH$PL��J�>�z��\_{�Lq�i��zK�䕋/S������xZf�G;�0�-����<25���Mi����Z�xN�s��	m��Xk�23���FYm_eZ)��e{[�,�Yg�sfZ��������qL-4i�׹��e�jߑ֊�R�2�Z.�ˆ�E���b�FYmk��X|��.	S�&�[d�Z&��jE(J�*#�MaF��Z�{�f�F��f�E�r��<4a���y��2ճ��ﮪ�]�i��4]w�?fZ#;�j,�e�׮Z)��e{[�,�3KM�Wj�Q�]��Xh�[V�l�����n�Qb"$�����
����p�Kk#;�VV���8��6����+4�G�����L�I�H�DhI�����9�/ƺ翮���-���V��!wuxZhׂ�צ-�ղ��E�a��k��a�8��h���R�.Gp���0̵l�ia�kqR�ˆZ�E���b�FYm_eZ)���g�2�eEh-
�#V���IA�H۔�-!�8֞8�s��a��m[E���3�xCZf�������ǆn�E4҂�R* f�Re���Ci{|��v�I����wRUۘ-�m��Ҷ���pCg5�3Җ�כv���٧�{���Q��F2����jy��Dm��ԭO,1�2�H�"��D�-Ωr�i�+t�{�����	��" @�	!H�b�L� z��݇q�lvr��[���{|0�^A��8|��l���08�ܶ�Β�5.�r�&6tCy;r���P��ˎVM0)���S�ơ�e�������\0��R��!��0Z9��SK��Ͱ5��p	�X��.�a(I�p�U~�=w.7PC�`죤�9��o��w��Y�J9@�����h��a�d7:�u�A�:��xU�MB����o/v:�PoWNf�h�:w2w^N[I2�a�l����Q����d�']�]�����bw*d����٦�r�S�l���x�u���ض�i��u=��e��s�����l�]�5��2]ذ7n�N����76�S�Y�]o<V1IE����(�m;y��]�vs��u�Ů����[��@P�8���c�e罓��d`W����f��{|����b�q����Z=����O,wFa�ٹ@[)��V��2����nꮥ�Y�z�3��"]Bye�ˤ6[Gu�Xf�k�w�[���u+�Xޱ=��h������3����#[/���Ǭ�mV����&4֞<��F37@[)��=�6��N7U�Е����γrT�3r�c@@�襺��[x^����S��X�kx�A�fYmr���OU�Wh�?�&�w�蓿�m��ߘ�se��6��=�:.�7R%�s����Q��ōW��/T�~݊4��Z��&��\�,���=���UHo�b��kG�v!���wnJ�u�3��V�����-�-�0+���,��=�f�S[�qWV��a�h~�������0)��ٛ��jіa�)���qXG���7</:F�qy�W^�ڱT*+L���\0��s[�#Fꎀ�3M��
]:l�U��`S7u�J-�kVf;�Q�}��#����쐩R;�,��t��hzͨ���ܵ�c�'׹�/+Z����*:�uNd�ռ�1���"�޸� �"=��Tk&�u���*���t���k:.8\.��̾�a���0��o�0)��� �8�t�)������n�(���F�,�
}I�P��=�F���208#����]EM�uQ5���v�6�y�7T$Pr�%�Km%��Ȓ�Q�a6���j�$�̰=�dev���ݷ�e3^�DC,�G;v�����p���oCYe����U���̴{޵�a��B�èL-�����i���ܭ�Ӻ�u�6���wކX��m^y@���g��{�/k�b>���{�؅��۹��tK��5���D<�͘]�N��:h�&�l���壌k��廷x2�6!��˔�h�.���7q-u��r�7l��u������(�kL�uu�.v�k9�/v��4����f9eVw~����� ���h�n�Ī�λ��r�]ae��n�6��:h�H����Q�Ͻ*�.Yu%� �L�w��#F��^�mF���y,����*���kt�b�I�<��!�ܸ!��ǅ�7�
��k��7�A�[����qɹ�����}�3|w{��N{�s�$��Ã���z~׷~�8x����)L�x'po���e2��Xy��X�Ú_�$8����̭b��	�m�J���ڭw�4+��"OO��\z�CY�R�7/��[q�T���ܨ�4��zxt`�-nN6I��kֻ\�[gb*h5b"�2:�9'�7�)M�7`��8�V�� oX�G���
5e�l-��3�R�+e+7h�����d�ui�g�%��f���\�����5�h�;Q�B΂�&�k��E���PϨ�z���O�˿Jw:3�cs�1w�����_����{���I�}AI��m�[��<g6�T�r�����lI���ʷz�IW\��4�Σuq�7]J��#V�L�_9��ۥ��������i4ҹC�P�&rd�������v��z[b��m]�e�yq�k�՘�Ȝ7<7:���Û�6�[<zuv�m�.�vx:���:���T^�(Zݑ���{�6{2��OX��g�6�`ĕ�C=!�f�x6�v���թ{{�T�X���]ۘ�"묥�W��r�9�ћr��]vton:���h��퍭w8ܙ;j�=N���\��OFx1�`��p�"��>y�=�+�y�[g �k0Ÿ{k�ͯ]���i��ͮ}�ۮ�Ű��h�1`J�L4��z��Od.xO\q����Z��s�۟\�-�0�S�on9�u�9F��k B�Wf�;;U��q��S�o:�a�ɦ̈v�R:���d����E����s�6�Z��yJN�5�K���<�ځ۵��as��}v�����\��9C�L獞'`� �c5�F�o��k�@�C�n[��.��Q�Oыq��,ø"\�\>w4t�ɧKnS�=׆�mG2nԍ�[v޺8�8��5�P��<p���N*;���\���X��-���N-;b�/I,��[k��	7L�/s�f1����JC������yml���q"�P���*TH����V�t���W<4���Y��@�=���~xQ���L`����B"���n�X��mI�mɚQ�[Z/@�-X�����OY5fM�vL/�9���9,�W�y�u���w]��������N���+R��m8'�rN�����12����(ǁ��l�O�o\$"���f���`�&����,)s�ɀe��kn�����28�[�X�׻������=����9�N&��ڑZ�bb�b`fQ�+S.vg=X����x5Fs����,O�&�qO&4�\)��T�A�]��t,�ɕxE
0H���3�/ɲa���	I/j�]`��r<%rݺ{\ż�1��HwUW>A����Aj�B;nh��U��r�Y$p)gnri�s��y�݂:�+b��'��H�X�7��G^�S�}u�n�r�ڋE�5QmF�a����XA3bc�
J���k0N=Mg�S��kvG6��6���Q�֮�6e��LR-��:�G
�L,�����M*gw�4n�����f�L
��g����`Cg�r�o@���Z���\ُ{��*Gx=E#�Hm-kV�Kݻ�t�5��hu�΋�"4S;�Z�F�C.�ˈ��o��ц��H���_czݞNKG�J"�	�T�-�hzluVJv��m�m�F�f���h��u	�4[^������,�r��!-��k����ڣ7|o�Ᏻ�Tt�vM!NL6+����,�/����bs]q�6U�q[)���m�Z5h��ƵE���Fi�)���f�0��KG�"��o���n,-4i�����L��FHxb���"0��sh��^�X�m�� �(��{kMh�e�4S4մ[6&��Z0�L��һWN�U�i�M^��F�~���Zh�ES�SE3ͬ4e�m/��r��i�k0�YDb�� 5ӹ[�d�49r�{��ƭ��&%�4S7�8��\��F�gw�>��uu���MN�Re�[7�Z�F=�h��n�g�5��u��U�a���R���Z��u��߆�Q0M8ԩ���T���nhm��-���T�Ed���ἥ��[Sɏ k���k~W��]o�x�8�E2c^�IW*U��5�)�-h�s����u�S�u���cOx\��t���"2����0��v��L�dxh���Z#E3bֽ��D-�˺����ݘ�u�yB\�e]IWn^V�m�����L֩F��U�\<�Xh�w{���4o|�un��<"�)��-a�	�Z7���L�<�a�ԴlX�[5Ώ�#�\xZh�EW��m�g6�ÂZ.�"�)�֭a���=Ue�+�\C-��,4F��Z#�06�^������i��Џ���fd�y'5��җM��+&�
92��}}r��X�5F�6�5�~X�*��S5���R�w���4W���O��o{���4o��)��(�;�c��KM��(�K%tqQ�ed��(�R�Z�5�<(�;��0�U��[E3�՝O-h�]Z)���k��7R.�Ѧ�����4[:մ[F3-���v���Z�˄��R���h�w���Ƃ���D�S=���]�[K���r7v�+-@ѾKٍ����n"�p��Z���/��]�a!�����)�Z�	�<"����̣Y�O_�5no8]UY�f닧���Ef�*���ע~�I^6�|�r��Y��VA�E&x����Ĕ�!���t�d
��]�6�i,Og��;W'�zو������r���ۇ�[�.�p��+�!�ף����eAu؝�;[�;g�<֎F�< g��ݪ�%T�7ODb1&�M�6 6��6���w�9���9V\�`m=�s<k�,��%��wR��a��~�E����񺳈u��
4>u�U*��iu�}�k�ٶ3-n����a�����%2��Mh�]Z)���j�q!�]Ţ4S9�Q�4g>&%H�wxF�&[\j4[EV�q�����[@¹���׽\��T��Z7�E��{��gR l�4m��,mވ�G���M*\D��޼rK6Ė���5�^1�z�k	�ń���WD�Gy@�c���Irܼ!{[�=�i�j38T��P'3���oq����[�ms��cu�y�z�]��m 6�i��C`6����HS����Ćs�Uݗ�*����owb����V���8��G
�ae��+���F�g5�4b�����Z�@�p��$&w���f���)#|֢ú��׍�m��C�u;q�cR�
[H��% ��u���%�kW�sgPW7pQ��խ�.XQ�|���A\�.��kLCäl�|Ƿ���M*���q�Ⱥy�_L=�o3��;�	�Ț��S�N^��9ռfd�:ڈyOW��^X��I�6$6$�s�7�ْj���)��6��h{ۙ�jۈJ!���� ���xz�`��v�&l�
�v�O\PO�E[ur�XhAh	��Y��l�{����{��풄ZGz3{�[y���Uc����	,��UJ��-����ge��`}�k�8����������'w���Tf�bk�o�Ȩ�*ؔ��N�nP���N��KYi&�@� ��)y��K����5���	3��D[���=8��\�Y�ɻy��Q��UP6S��ۧsd�4
T1	����~�]�SKZ�sپ횽��(�×��r�Ӓa��;j> �\wb�{Z�#GyH���}��T����#��3�Z]���D[K���g=�UV����g��J0����R����s�Du�������d�-��+a�+�a�{t!��́%zcg.]����]���ɾP�L^VYzz���=u&}u-*�e!9�{�s�dCBd�PH'/��u������خ9�Zk��{nwb���nk-��x�v������Y���Ŭ@]���{s���m��)�7���L�����Ĝ]-�1յ��sv�p����YbG�b1��.ݕ)�6 �u��{&*�,�b�Lx[��%��ioԭ��3 ����� b�Gk����{��˅J��X��K�4��֬���-��R�m_�[.8\�S	��Ѻ��-���XbyV!����.:���� ��s�����[�fD@�[�������ԫ�"�^�-FD2�ʰ~��g�m-����֩ZZI�89h�@[FL ��
:R���G�m�/��ٝ�����Hj4��Z�Gk\�F!(��2<"ۨc��~Y'n���F��@t���j�9 ��f�Dq7�wz�s�#I6%�k�R-��R�#�̈��"��sݺ�.�.��z��is\�u!��ʱ�����׽�T��-�$0�iF#yԂ9�����p�Q���^$�wWw������G9�l^��wW`3`t�]�T[^j�ժ�v(]�w�������.U�uڦ�Z5Z�0�{^��
k|���:�V䫕*��ݢ�A���m{:��Fwv��T}��r\܊����`t�l�\*]�K����z����oo@<2�G{`�ϣŞH�g�����y^]�W������9�z���2�/B�~ܞ�¯&�RU��b�y�<��Ed������br�w�˝0�eG0�P˄b�$�^fM�݄�sNu�r�zf���W��H{�[�玃p����lf�/��LTvu�f��5/_:����	E����4�.y޸�
]r�K�Z��7x�U�0.o�6vj 2�T�7�w�A�&bʨ�Z��	
���p+����VK�iǱO,Z%.NM��K��G���w�|t�f^%W@���l�˓9S{�Ry�D��"霑1e.����;��������\�|�����5���M��~v���|x����O5(���[�2�*(�{��\
�h{{mB��>�Ӭ��������S����\��D\��]q08�"�mq,�����3CՎ�
.@̪錜�nϱ��"^u�Y�Ŀ�Ho�=����1L��C�;�l:�L!q�M���>�q�1t(3�#9h2w�<}:�ӮK���/f��P{�}#�<��zصRO6>�c�I��]Y����p���&	�;*��;)/�l�=E�J;˺��°l�3��0b峭�2ӣ7�<D�}���w%��"��|R��������$�a@hMN#�ph�ˆ*L��\�6LU�:kZlk[F��IB5���"C�)z 0}4����H�knfy��0����F���Ѥ�ڎbu?�_]s;���6�b-��{^�z�^7�}��ig3[��.0�������%����6��{��8^�3Z)��uV�.�	e�g��F�^\���-e�x�&���0���h��V$FV!�MݞytQۖ�s郎�����I�7�?za��5�a�Mn��LQ�gw�F�F���d�`�Yi{��~��o$2і���ZQ���ClK����H9R;�YiS]�JڦkZ��C�G�F�.�XF�5��V�Kp�n�Z [�-�מq�}y/�G�ӵJ5b��MC�ܖHژ�Si�	�oaʀ���:�d�Y�Y��T�=.&�)B�� Dx�]򚤭�ek�ܸ��]˼"5����b��b�T׵�D��3\���h��ӽ�1&G܄�QZ;jpb(�HE XKt��<c��$XiS[�Jڦ{Z���ϻdj3��_$wWN�r�k��"��l7�hny�����c��o��V8�K-S;�Dj4ktF��L]�-a�M{[�KS+]�j���%RY�G�ކZ�.���*kwI[8�v�j���C��UR�Z�.�Z�*~�ky�e�f�ڷ�ְ���Db�4>���N��6N�<�]��'�b���u�{I�������[�n\�c:�:��e��ط�y��i�v���C�^svZ�۹y�g۵�9�.Ƭtn�B����o���D���kp�p��l���c�Z��ƻnc<���m��F��]�oQ<��@���m������������ݣ����eG���t=P.*��~�7��޶����-���Q�Xis��iSZ���u�\���Yj��������j4��b,4���#�25lΧ�n]\�xF�G�Dj4��j0�[^���T��!�m�h�˒�I0e���þ�b�J���V�5��j٤��(�Xig�ݺ�RI���5��,5O�3r�r�[�wݻ�9�����$1X��t�hUVAG8�eB����� ���mw�+klީ��z�ee��܂3�.W�� 
��^�c'�L��D�S�1�9�)@���[�q�t�����ǂ����z���hM��ƚ]�ڌF�v!�9�y$�h��9�Y,�F\�+b5��-�aLרhzբ�S~ת8T��e��:��Z\m�������b�qk*k���9.[����3}���k���9|�2�i{|�XiS�3�-��5�6aF���V�T��阌vs;G4��+(���F���3��:#5��6���ԸU\�*�Z�/{؋�LV�{�ҍS7�Dk��j�lR\���GwuD)�,���s��a�f��ٓ��w^����_����ĩ��;bg^FU�Zo8E�i�-�v\��o]�q��I��Z;Y���4����;��Ҧ�|��AՎ��Y~Be���a�ѮQ�.��������l����V]Kx-��"ؼ���ykLG�Yim�f�H�F��]�:q�u��r��A�{�2u=�˻w*�U��Q��KQ�Mo:�KS-���2T���O7$�����������Ѯ��.vZ��+kSǩ�	.��	e�aˤ6��U�CG�����E��5��ҍS3��ܕr��#g�R9�0�[�T׳�D��o�~߉���g��㾴;jf]��hh*��q�e8�a�{F�ww�f����tD{ɱ���g��b�ڶ�Y�˕r�I0fR^�1��pLS7�Dj4g�F��s�q���E�aXX�)K`���sV
�l��]U��������%����Cj�=Z�<ia��sa�Mo}:�]V\�0�Z�s��4ktF�K���J�ǵ���̵l�z�Y#���!���W}5[��uST��w��ot��h�Ό�e�Ƀ-e�$4wص��5�o,5L5t�ճi5��ᖣJ��U��J����J��aiJ�Fcw�Ï{y�8��z�U���?J�.ُ��v3r#�^9�\c/v=Wgz�>�E��L�^�Z�* d(]2	��@���#��c�f�ǫ�Š΋۞Ck�i8��Vw�s�������W>;n��^ܻ��N�@��z����W.�v���@�[̹�64uz�흱m�:Qt���{��Ë{�{��z��>�r�F����-��������Ӯ[���T�]!�m��j4��� �ZV׼+����zR�B��x�������9�Q�Mg��4і��t��T�G�f&���A2*<���,I�C���V��b3�}x�A�g��{>X��k�%�[ �}�1�9sq,s�pw'=v����Vטzr�/(\��]K5�.��{f�V9��E�dfG�5�m�ؾ��7i؋��+~K�u��R�\��4��e�d�}�>�=��o�t�,'�6p��y�+\�1;k�hH��=��<�q
w��u0�I)��U,��ԢO0�6�+�e������u�ȫ|q��+3�[�c|�l۪�,5���G��C
�/gQ�HFj,��癷BR�SW�Nr��{�k��\�-2����v=��� ��ƾ�����P��r�1�S�TȀ�nuD�Y+�*��CnY��Y�3�n�H���p<"<:
y;�[P��� ���bG����ú"�A��{R�����z������v)\UZ�B��CҗHpm�;q�SF"�}o��(����7����Ja�a'�<�df5���v- 3�cM�M%4=�g,�>��\|5l9������J����b����EV��9��b{Joo{���=��p4LL�z�eA�4���$���j?3����mFe�|>X]�g�|.�k�7���*�h���-��3����E5(����҅Tosuiu���[qy�JfOFk�yݵA��xL���*_rQsO���[�u�4q0ZE)��yv��W�f7tq��h��>���i͕�cp��0��kudm�f��-s+I����͊�*<��@��3��Ι�30ܻj*����6Ȼ���h���ijb�o	�;ȉ}x�n(�V6�o�����ouHW>$Z�>Os�=���lT�<��*?w�9�76]�ܷ9c/��1y.'wgo2;���Bn�yQֵH�5��g��f5R�.�3�%�y�8)���E+�{��L�J�sV 9	�.���]E[ޥ���w���/\���\.�=�V�ůq�߼�N��.x�3�;#�;�nk�H�ZyH�v�{��gx�*��ʴm�2�j�p8 WTs��w�U(�ꉢ��P��c��[ڼv{L�s}�\TJ����1Ss�X���"��=�J~�Q�p;[qq���Od��#p�2�0����J�����Aw���wK���,s<�� Q����ʄxx�+�9՜ƁѣϓPcybV��:��[��:#���F��y5ڕ��Nٹ3�M��s����.-���smVR0vYH�e���n6�z�;�;�׃)���m��Yͻnx����Lj[pq�˱�uvm�&�M�6�p�����q�s=�a�i7I;��F��N������P�G��������8fz�e�����l]8�ktGc:��n<�r]]:۵FSæ���c[�����Z�'��$�8��{�3���������M����.����r�z��&3@Y�|��%::_Cd��U�n�4��ćo=g�En��=�.�J�]m������z�#e��������u���ݬpv��f�M]��ܦ3��')�7&���\���V��_#�1́!)����u5��-����731�vŭ2X@s�l�Hn��]��:s,��j*���d���>,��"��M����V�ۯC��m܎��l�s�ܻl	�,������=]zL�	uvιE8���T��:N3ɰ��]sV{<N�궵90<�*�$4������E��B+��|���S\>N�D}2�9���qR�D�&nȚ����+�6b��n"�F �<�2u�@u�\3�=Ձ��-�K�*�@l�	���z��I$0��U,g�s�>�v���ʉ$B>E!��°d	���s_�|�2�t �;:�VrnoEtw�^�]���SC� <є���v�r��|�)�[[3����.˺X:PM�s�]w��n�,�f0;��<�{S ������������v.�O���j+���� B,���JZm��������	@1�5BMgD�ŧu4�7Z�D��w&V�_`��k��?��nt�E2�sY��v�$q��35x���"�BBX~8�D�>pc�W%)���3e9��2%�:��
�'�#��)�������Y��1.��qֻW�{<��Ϝ�o���0�P�n�n4��tF�ح��ثj��v���:�Id0ca��kgk�@��ַ.��ˀ����JF�G!mV�ě�i�4�J4���7��o^
Y֩�`�#v�E$�,�nс)	a�ǧI�Z�΋p�*���YMAi�������U�:��	��6�75��q���^J�J�֌�(��D����uiu�� �\���S�Q�Oc�����Gw#���I�-�|x>u�hN�wd2t�yĬ(��m�Uν�'5���^���ָ��S0�n����@���X�ç`��=�w����.����Qs��(��٨1{3�7��.�@�UR��_Z\<~���e�4�+��y��pyU}�����
[s�.xpq�m߼����p�j*W^7 �����SY��V����%*����r��B@/*��jU�3�����5}�p�=n#3N�P�11ۻ��9)ģ���$��o��ZDOF�sM���9�p��_Jx��q,�����2	�(M**�2�����vD�ɬr�U� �59�޽�0��m�wx��n2���A`���]|���i�;PQ�fd��[iF���3� �[0�|=l��OQѝr5��$2�)*���#�O}'1o�)�Qsz�y�5V�V,��`,����vkq���z���Pۜ����qx���fl��.z'A�a|VS������T={QF�^%8���.v�D����#�`�Z�_vu���9$0��I�7�;�̬wR<$g\8�-��S�ʢ8m��IZ��5f׳(�@�����?E�aU=���[dg
��. ˗�-����Wf��(M�SG��x�M�[�F�e0�0�� �⭭�o<�a�َ�[L�9�g�۳1Sm�ܲ�q���Dܖ��G�b��M9t��y��=U�cW<y>:+!�����[��5��*	���Y�{=��H/]y<p��5@E�[eh����Y������Df��pF�]s�ZE��{Bk�W��N��H�%�Q.�.��v��t�wJq>��u�����:��։ЎX�.ڲ���ct�)��<��%�@�;H���h��]�R�`]�%����9U�o�g7�i�X�I6ɇ1]�@oP]�u[s����ӧ[�(C�������O[qY���-"'}��zV�7�k�x�d��84��ڔp��.f/P[m`��ߞz4�-�b��(�TPD��oVGIc�I 2�n��U{��[��$�p�Ye����y�`�:υ�3����[h]�/#ao��[��k�{�����oY�1{�qGMcm�b3�"��%��kq����6~8�L���7v�x=r}����e5���f���
>�y�^��FÄ�6��� U���kuskk���P�1�Q	`@\zn5��L�f�aK�����{��l���rN 6�{�o%�j
:���DE���A�q
�v�/��"����8�ژ��:�h\�;��{�9@�~��&m�EU�z��H�bM.4��l^hf��L��)�=��XP�-O�x��(�ʙ:���{X��%�1z��Z�=x��- ]�}���8��"�<�gXJ:0��������g�w7�.�Í�(��Rz�;�(���V{��X�M�ه2o�\]!����9'���Í�!�bt{ǻ�ޥ֔m@�ݾN�(uY=ʲ�U�Rf򳍍AѺ	�Ɩ-�U�+n���U} ���l ��b��;+���-Ʌ.�������ɘ�W��X��%C��A��0�uך.�lX-u���f	A��K���';}�r/��Anh��#����]�ӔpxOb�0ᤐ��1Q��Ws�}.��6S,�8 ���U�]+o������7
O^7<3Xqٍ֥V����&�tƉ��F���Vӆ��S�e�=F��g���L9sR�=���ry�(�	���jES�KpW�N�5����m�yϝ[w=]r�'v1[]�"Nˍ����D��pm���R�gO��NF��o쓞�]���g����..��z�	�ε�:9����ȝ���F�mmii��ɗ]s�i���۞�[�3z۪+l-����׮��U�����W^7z4AH�4��n�7�v%�����eiN 6�y��oG��aGf7#z"2�QgG����w&���Y'OԚ��jc��32f�-��=�����n(�y�E�wi�\p�%aaD�B�O���{kgp. �PQۮ�[M%7�ë��ɋ�"f���'j�E8.�5G{3���N�����K�]��.�����gٍ�����I��c�վc�=ks�<
����,4e���f!��g���R�6�- ����r=����9����o<����3Lok|�}�GM7 �y��Ԇ����̓rX�z��Tp`ܱ��-adZ�m3k��<���8��ZJ_j]�Uˏ��wi�5�-�pL�|���z��3xMM�ݞ�n���5�<Ϲ�R3�ۃ��t� ���}�q>�������B;�pf�z����O&��7�`�8�-nq��y���Z��N`�s�~��~j��j��O�*��Oc��v��9�SZT凷���{dI�z�b��n#5.��g��^Z]�}��;����3�|$��1u�d����j؊G��ܕp�]�nW9��"��w����9ApUF�5�	i)��^�twEmTó�2&1ļmz\E�͋�Ժ:�jo^�$�����g5�p��hc�
�奔�Y������Uw��vOO��o3�Aи�~h~=�>2���y���8_D��&���O[3Ggip����|�b�	g��V�\B�	j��
4\Υ1g)n�����uj8�܎y�c{I\���8���&Ys �9��5(b{p%�	����S����a֬�&�Ɲ#&�tʟۏ�/�{�K ��E��h �?UX`y)EF{�1�8��ٺ��Ps�sF�,2檅/ t�
��)K�x�+������C'�.a-�	;��y&q��}��@�o��Y��ǌc(�����߱G�����5M�ba�XD�Q@N�̫����
#d����]KIAI ���@��,�L�5fNH�f��f7��C���h0��3��w �f�i���k�kM>;�;���8�X�aEٍ��&�go̽Dnz����B�;z���*�1'��z*��Z�3�C�|�%���B4�ȱ>g�u��w5�1�<�r��̛�-��a[���K����$��; *�˶�s����u���u��ք؆и��lIS<b�y��x��j�J�v�� sXWi9J��u�Y����(��9oR�8��=r��W�m��8�mdݟl�%ٸ�ݮۮ6B���SPR��J,Z
7���Ԫ��Pۘ�Ǡ	7�.�ni+�5X2 �B4&7y���xv7ד1C��p�@L6'��wL�[q؂0��u�6Z�0#U���{3z,ȑzvS[7]<���,���>s�=s�~+E�^��TV_|��	ߓD9��(�e\�|3�fR���|��x�XJT� ���+�
X��*;4��U�[w�������(�Ze�שa���(�C<���8M�R�Ԯ���=r��R\	E������ģk���zS|�@3/^�>�o�=�uk�'� ��Q�zLQ����p���:�Zf��P��}�ViE�)�{際�B;���g�݅��եb�d[n��Y(�M�2A�+Χ1.���"j�Żu�ם��2DU+��M���l$�:<Y�c�c$v%-��9{7�t�X����b�z룵AZR���9U�ac�	?�maH�1u�B�ATP+n�5�v�����S�׏,��D+���f�'k�y��n>9�ɐ�6����ޚ���J6����IK�J��&���3}��p\4 =�F^7Z����/��-$�/�[������v�a-]>�,��U�Q1�\U8l�ع�W�XD��!��n'�I�A;�Ae5*�Ę��j�Y�y�^EOER��u^��{�Syډ�H�T�a��fwsx��TU�}0<)��M0�Sz�m���U��{�E(i�_��}x�	�6j�D�Y�)�� �^�N�]ʶ�'	��c��	��8���u�G�D/?8�\E�f�@*��(��M��D:���7o@��L�lt�	B3��7��9�;K��Չ�[%'1�!][w�}}f���$��^r�SSx`VѾ���˫]�x7zTL�ӥ9���z�v�u��Q�F&�l�6���wnҎp�)%<=��f�n�Ő�ݥ��Xh˻J3��cq��֥�©�4x�:�6��uz�.�_hQPN:R�-(�i��ɶ����z�M�9���*!�'�����O�}����0�B���5'}��YiE��K ��9hN�Ct_\�L-{�h�z�@��]�u)�r.�,�<��E9��<�53�ng���FX�M��Ѽ��=�8�������]��7m`���y/8�%E�74a([b�qt�e�Ye��G�y��ƾ�| �ڔQ����*
NoV�3�TO[qY���}��ܮ�n3�3ٍޥu[����٪�e��]mg��ɘ��1"���\=�4:�� \o
�]mEP�݈a\ӛ9 ����a=�����:Y�D�ir{/��o�|���\V�"',%NW�͈G�pv|�+Nێn����������r��d{>��n݇X6x�έ����si.�s�=R)�Zű2uJw���w^�J����.L�n�<���J4���<c93WV���.�u�7s��k%m^���(�,;��M�.�����Y�q,k��.�\<3-�ӱ5~�[���L��"��ΰ�YQ���N �JNpx氲/�� wZ����6RJl���޶�,�Ϯ�"bP��R���X���V	��@�RX"[��t9Tu�{�f��6���i�I��ƺ�B���/u,@{�׹�����&{�m��6'�0oA]W�*�'�W9�H���DD{��S�w�u�y��k�lA8�1�stN�0���v7[z�A	�Ү��Һ���x�%�Z�ڕ�q�z��b�o^�^c����V4H��KZq(m=sÊ�Y�~�����o��nQ�p,��*b�G�ȼk��Š3F�
i2�.p��)�85C�~�@~v��<8�%��o�{�A��7[�#V"�N���|	= ���IT��)�-�[��dLn�]��S9�%(M����|>�g��k��5:��Ӓ�J����U��(���c�M�8[�~����#����u�1i�ـPnz3_x�2\v�g���kz����E�< I�Kb��P��i�: ��̋n�zEF:�O1^�!͇+6�S|;���z{�oXQ�2���,���>� /��os�m���)9�Ի�a���cq�Z���_c���N�G[v���U����sD��_��7����z=&�)�FbL��+��x������6���i�I����h����}��D�F6"
�qw�=�.�$z��x���M+��k��ɘ���O��]��ٵ~��"J?� L�� ��HB ���*_���~��)�+�B����j�l�ěI6���ڍ���ѭ�m���X�h�U&����5[��ʪ�zͶ�Sj6����j-b�^��uU��J��E���77FBe0]NQ5�T[[[%[mbڶ�KU�6�U�m���m�Um�Q[Uɶ��mUImRU�E���mki*��ۓk[u�ήh�nusnMA�S"�isr�&��M�{��~-�Fo��������m�mV�B#��-�*���c��_�.���|?���!�fl_ۥ쯥h����5!եs:HB ���p���������	!	 h���%A�?jk�?�����L�	������	!}_o�?"w��#����>B>�|�p��|�2 �_b_�{EP�x��}Q��Q0
��gSI���(������߿��!!kI ��բ��-Z���F���khիQUmb֪6ձ�U����Q�mX���m���b�[EV�Z�6�[Q�cV5��)��ն�k���m�n��6��bM�����TNޓ;O�a��<����B��	!4�����~Ϥ��/�?�	���|��ب_a���$-��� �����B��*��G/��/ڃ�Lj�(�J�������X>�_�X��1�|�?p}k���a�I%������_Z�����k������?�&�����~	B@�?#�К"�/�|�!��p\B��g�����E �(>�����1��x�%��I!  ��|�K��AX��7e'I$/߁,pX�a��WaA�[�!H�O��~����$��/���}>�!/��][�~?U&���(%�~���>k���k���aG����>f�!H�B��l�:���B��0$�����4sB���P �h?ĤR�c������ϯ����#���=e`�R��/�A��_�Q���a�u�0/�[=_HH4�$~#��J���?������CI!	 �T/�/�Zb_!$+3�o ���>��P(I
Ϲ}ʒ�]k4��Ƣ�3�1/Ń_�p���?����������ܑN$�M�@