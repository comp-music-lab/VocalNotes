BZh91AY&SY��(� �_�py����������`��         8HJ�@_YQ ��!sϠ
       ��JP'}/���{h���;�E\��$�*��s�2��8�T%RW��׺1UD�|��T�q�D���T$QnnQO!-�k�Q�VtIJ.,��(���������QOy랉$��ܢ�
�t�(��h��<�:QJz����3�n<�(��#EQ�c�������w�tP
9�tQ"�$.�Q{Ց]��EQ��J(��Ί=E2�[����(��	��)�       S�R�i�F�1�4ɦ���~&$�J� ɂ�da4ɠ =��Ui@� 4�  ��PL�R�&L�41 L�LMO�JHUO�A�14  4��  BF� I��24#�L�m�z��'�pc��G.����4�dA
?��A ����UD���DA�����zO�+�#\�P@#Q?Kl�J�����(��"��e*.�������nH� "����fX+�E�Rx���3���'��ybp�����}-,���у���otJ�c�f0.���G��(k�ъX�������ʜ<-���Y^9b�U��:��A���p��1�aQ,k4K�9m撗F�Ÿ��	��S�n ���|p�ڍ�9��\2�+� x�xe���ie��䫌��2K��V��
޸L{�:��gv�<�[y=�ƃݩ�ٺ��ݝob�\<wF���s�6G<\wDRaI��ʵs\V�5)�s�W�W|�l\Ww��4� ����8N��q<4s��OB�'L�ۻ�7�'+��V\jL�t�i���ޅD�ɶ�Pw�t�����/@0A�s@v	ا6��L2X
���Y��|��2����!훃M��z�`����^湏tǜP��\�(֏�T�aߥ9uكl�)��u>��އon0��/Ԍĸ=�9m#q�&��a�5xm1P�\�w�6� MɷJ#=��.0�H7{
:͙�ub ��}5G+}�8h�P�eg#�a_szR�^}N��3;0n� qǃ �ʇM����|^no+8��v+:a�����@�f�pX�\P,K�*�A���U3���l\N�Vt@[BׅKRM��K��+��4�k"��ݱ��J��`$Mݻݮ|���
b�ii:{����$��k{�S��<���gs�W�����fl�;�I;���se4	��h���6��{4]x�EOpxf�x7�r[�=��8���õ)�EZpdm9nK�@�@h\�:�ծf��ݸd�wbY���pGt�`Yzs�ʣT�7��q�"�FNH�2�^�o;���;���x�;�sl���[+L+=�Y2��lK�6��Ih�d<�u�ոn��KݜI��<����x*����ټ�UډR0_���Hz�wD�w6G8$��R��Ĭ칽���Mt}��	�e����7��)��.�;���}����]�v]�N7�#��ab}6Wt��ȱ�>���1��'@���#��緃� �63U�A��ci�	]�t�ܗtv���x���{���p�y�/ rЙ��MP)�wv�Uv�"oh�8e^�4vb��ݼ[�D]�ܗ��r�wL,s�2���I���` &�T���i�z�kw��G\��� ��7����ۄ-S��}�oMs���Hҹ��L�K���*��+^�l�6�0��͡m�SE��[6����$�kEs{:�0�Ư�1���m�y8S�¹�ls�g	ϖ�<�N}�>��N�t醲�gf������w�-hф���p�a֨"�--$.�]X�A7%x�'�7z&k�G�p�nH�̩�⻳S)nN�v�3�ex��G����,�y�ޡ����A�Qۨ	8�o�Y��'+�^��D�eC�.�z�{�<�\b��I�^׶;V�q�U�ܗgw4pt�G�*��3�W#K�Ă";�{��6��V��Ed�#��8i��.�����GA34X8�D�����͍�b��H�秜�oN�t�d`;��k��"GwBI�u��k��c_B8d�n��b����Nlvڠ�q���6z�yP�ķ�p�cY��M;�!Ϝ<T��2�5��|7�$�Je�^�a㒐3['!Z3��W�v��s�˫�&�sێV��l:��v�\u�p������K������ n�:֞v��rr��+�:[�U�r��ॗ!,��_&	n�k�����ۨ���d�qM�z��n#Nf�7k�N<Y���"�fe�(r��w�rܠ�qNN��q<�v��Ea��=y��2��=�2���� @���E�7G۪�������S��~ҥu���ssY�a��1��.�<}7�G�q:���3S"o�u*�{�����'��sq��s�ؖ�<f^��rkXI�y�nq�P�t��h�����p�s½��mWkv<��ptg�2�oO&��ù�;�ˣV�Qq7/�co[s]E��c�&�¦�`E�5Д�5�6���ڠp�s�Ӝ�Xݎ�5\��Q��Q݅.�0�$1We�LL�`�khh�]��F�<b�	s,@jA�˰k
b�SCp�Xs(�q��c5Esai�	cI��v�푰��l�֎�n+z�]�=�k���99h���iH%��ɦb���ĕ�`����S\�Y�n.��Gls�W���8�-ɇs���Θy���Mtdq�ݢ+ؗ��x�'����{f�Gf48�U�;=YN�����n=ek���M/zE��4Myk�vse�^Mh����$V�$��nAơ��n��8�֫:�U5�a��ĵ���
 ơ��.�n�ٺFê�����+�b�k��=�:��p$tα���"��5���q�l2��qs���G=�gJ]�Wh�kLu�-rm�޷<'����/D�������p�J5gY��?g�����=��N�#�=Q�iGYy\m�n��t�<�d݀g��xk8wOU��&=8L:�k�)�D��2൦�ڄ�`�*�C2�3vG2��@��a��K�WU�@V=��R�ٴ=a��i�v۩��G�F�$6e��A�,؎ ͳL��Fl�i�tڻM5HVR:�J݀pu)au6�i tk�6چ�ц�Sz޶ ӎx!ۆ��蝜���q��1�n����\aC^u���n6����h���>�]�����5[1�)���I��SJ��P��	�r������W-�s�ƻV����=�uu���u����X�nW�W�c�(Ä�j[�P�԰�����X�
i�6��[3v4F��,
Mn�suX��q��)��͗m,ED�i�p�`ks����!n����
�HDH����k���Ee�
�Єˡ�M.��.3�6A�����鑰Y�$#��e��[��i�[=ў�j�ں�ycH��m˝�s�x�d@��W]�7���3���<�;v���eN��=z9&��s=���q6̴&Q�M\�eM���Rx9X�G��p��gWOS�u�8`��:{�]g�Ɖ6�rv���^�ڷ�CaR3,�w-sDB6�\mcۓ�V&㮯\�a.�5&�K�E��IKu�CmQ���+�a;c�=\v��r	�j��.�"��b����M\д����j������hqHAB��l�4 �p
Y�k��s:����7m����n��mg�5�抨�%x�j��ݚ)�9�p"]����#�rS��Yi�>؂Ɂ�B�ZlL�r������T~�AT�@U ���3��u��O�-��@��W	8��U+.�Z���?Q�a��^���ٷv��d��:�/w,�����S�1��6��K��o<���3Rw��� ,�9w,�Uj�''i�w;�>���1���&���G�Nҋ�?,ت��+��8�����I��&����Wc�=��n��7Uy���=��;�8�cg��]��{s�kyza������`�$���f�F'���}f��d;��z�'��!������<�(A��h��0�n5�����F= ��XH̻��<VڳD
�^S!���쾾ҝ|�*.���Xd-Q����S�<f_�\���]�/o{fw="����z�~]�v{�f^yۗ��*���.��4(�lI�{�����h���<��;gM}��ɎO8�~��O8к>�-����=�!���e�q�.GA��np�� ����;������1����˯�b���=��:�i��9��˾>��\�U���������k�ȎkZ�1�h"��#G�z�����}D/�_�wL�`柟�7/�؉|r�v=�r�S��rtk��產
����?�sF[z�wݽ��6���Me~�+]��U��n��فr�yN̞��wǡ��Z�f�;��Ο-������2�ü��2��&[�o|	�'��p;@*ft�߷۶gL�{�j�<��e���`�7������";�w���~���Fݝ�0�ɀÐ�q^u��ٿn=�Mt\�\ͯ�!�Tv�-��}���w�4^ó�q�������jvr{���&�t��}�۞O=��7�r>9I���e��B��/��{˲��8r!����ԥQ��ݓQ�K0e|gݫ���A8�%=�>]�-Zb�3�+#�y�T^/��t��/mE����Q�Bw�Q�������.N<�<��E���:�=
�3�S_�޿E�����U��v(f�rő=���}�Y��WE�ѵ����9��o�`͉����ҔӜ�]���a�������^{+�g���[�G��;�x[�-��	w��� �]ٛ������l�|��9n�x�r8��c�;E<g.]�;��֥���^�;�@��)�-�R��t������ӭ�qq΅�{_y�C T��������C���Y;��ٓ"8�{Xj��A�=r�L���>2|Ȓ���#�qtNM���z��=��ӳt���j�:�����`���w����}旰��e�~&-�?a3�^~�H��I��e#@�G2Wn���ېb�f[��{�����̣��t�������qkk��w�C	/��{"��L��fh���^m����;��;=��뇣�/��>�<GY)+����:}���ݪo��B&��f`�}���uho�w<H��r�]��$����vG�+z���Y0�?iFwGǎ��랐�b����:�8�ɇ�^��A�v���j�|��V��k�@}	�u�ޝ�^�S���o3�=��?�4�~�ٙ�L��<�ex6��OQg�M�o�A�ֿmvu�{	B�}*+����uou���_$��� �w^u��f�u�]�}�K?0`>���;J�>�=0��s��<:nl��F=���9�vk�ԡܯ��*�}�s�~� [�$M�n#.@r秵�/nv��7Ƃz��h3t�S{���	�m�����"�5?S�@9���޹���W�����Θg-d�Nȼ���Pe�˝8���B(�������ְ/��ѿ{��yЇ�%V|U��<	{=y��2(�\F��h�����Ę�^�E�d��7�Opݔ��Ӟ{ց��Vʄc�܊�����y�l\�x�1�8�#����7Ἴ��zv�y��}�k G�"�{�^��gXM*�����5�2�g�'��@rEA ���`zcx�����P�V=N|ߐ?2t[^��C\uR�y�ݔ��[y�r�5A�=�)�Oli�-�X1���L]�!�fgMb�Лm����6�;�8�'h�������:1��m�,T5vҨsjH��2J��Mr(V�nއ[��u�n\��T�m���$������K4IfAQi[�CM�:s�^���=]�qX�΂�٧�׭얺�%=�1�8L�9g��������ǎw����Lf�ϰg=o '#1Ҭ�������o<�;�|�x�MG6�]V`�_';>��Y@�i=��|�>���>�rz�7�r%
w,xkg�/�px)Ĭ���A�<Y�ӝmͺrf��挷�����r�<�4�]Elro���m��H�2"��B&W�r �g�A�x�1�M��իW(�V�襎(�hk�KFx�Y��n6*����"ZV� [Nin͇J4`����z��D�(���٨�T��ȹy'�l��3��1���-�K�s�6 �d�Ύ^�۝�Bj�6�Gv�Ywa�/��lhW��de��QdK[��Y�zf�� �a�3�Kk�k={wd3S�����ݳI���az� �{�NE�:�#���-�l���K;k7���"h��䳿-AL��O/X�| 5�ee��sA�Q��Z�[zk�gk�{��q�]D��X����Y;3�l�����T�B'��d#I��x��Lip�aI�T�L�1@�L�9��yVjþ�g̏V����A�u���\�-$��Zաmr��
��J�6�6�@��ͻS�9���@V�mܛ݉�dUm����)�b���N}N�%U᪱ϻ�і�U�D�LX���������;���f�A͟{6��2Tz�K	�����5)����ML�볘�\9��֣����p	vme�>��=u�Ia�8��ҍi�1cT�"r�
�/A��gt읯]�7a�OwϏ|>/ʸJz�y�
�ċ�z��s����K�����q��&�X��x�p;�|ʁ�g�ܸvbr��B�9\��y������}���m��^��{�U�{(���%X'�~�˸�{Ǡf��ų�0���ݖkv��Z��]c�?tԅR����$lr���ݐ��x!$^�ve~	��.<�ʄ����a����H����fq�$Dh�qS��
`QĘ�J*�kH���4hC\��=5q��������\U	-`�A��d�7�4�53[4�0�q�9��xD�x6�8�m#������2�]޼Ͷd�ܖ��/�m�)��d*��/^��өC�LO���Tb"7|Y�0w�b3/�j;v�@�X�0_͍�霌��{jT� 0F �,;6�^ F)pl52|���Ӻ��wC���g}Ok(��q���$�0��M뛷-{��;�9�;E18K\m]3�Jkv��_>n*������@[�Bٹ~���+�!ƥ�Zr�[fW�L�y`��ޙ;����Aox�m*veQ�����CH�Ru�(`��{W����th�:A�x������f���N���r�Cn*�^�0�!	}��cU�b>b�y��lZf�i"G�b9��p��f�}Q݋絇���L+ύN�*����&Z0��_1�����_i�ǧ�d�,�a|�s�D�����s�Q	_�<1~�-Y�KE��c=��$MZv3<x]��|�]�uy:ty\���S�z���Gb9��׊�~�r��Fe�=]����b�q{��K���nn���A&0"��=��
��
��gN�Б��&T�;��3�Hvyf{p��NM�3�Tx}۹���`o�'ޞ�|䪴�*�k�Ҍ������nsTҴ���8́_xo��{�::p^{�ۜm�C�c��i��fa��	�9�oIC����Z'����zB�r��1 1b�b�7�gfT�~� �U��Aq���}�9��'���b�5�	�����f��'}�����
�N�:��k5J��C�2�?G�
L@��H�&D�S�FQF?�Ă
�]X>�"H�|�nc8�_<#G�A.!�w�@A�X�I^55�s<㱔�(����X�$�~�t�4�g��^V�X���-�2[mw[
j�#i#"o�Z^��9E&�@�T1�!h;D��P��v�L�Y^Յ$7�TL�F�I��$5�}+;�Մ`!����ϑڐ�>�����+V�4�3R��6d�n��16��<7�T\m6���P�Q����uޤ�����]�}s��P2b�:����)�R�9�j��`�k�M��e$5֓5���*x�Ψp�j�2�%���Tx� �o)I��-|oW���^��h�uJHm�a�&q- ���o{��)7���4Ґ��TѨ��I�6���pE��V�؆�d-�yI�b�43�D���~��;����n70�{hFO�MɎ��pӎ�o=�63:�����E!s���x�mI��;����XRGx�A�RTXk -��RC|p�U�� �h��E6�C8�X+h���m���F�����T6ڀ�M"T�1���(�1W{P�9@*$ޒ�a ���_z��U�0$��R#�2�h��@Ϊ)-|����)�+��(��"怇�D�P����V�Ouc1x���B�gd0�[����3�Ɇl�v͝U���t��M���s��,�fO^Z�| �+�P��k2ٝ��XG������^TQ��V��d�C���rF�0=1ݤ�QXQ�^%�5�a$�L�GzL;����{�m.��"5+� {�.H�+{� ��4�,w�.+f�uFM� �b�,s8����xw����#�	i����¹#�@X�zy'�Q)_���a��3�U���:�U����U)�,K�w��=�G�aGC�S�f_N/ Ɨ��h�,���d�L����=��W��Y�X�X��"S�z͇�����f0b����{���v�Xv�ğ����Dp2�w}!7�(TЬ���IRX�+��dz	�,(���d����FR<Q�i�����-�⒄�x�x�Aot�;�� ���\Q�f~,5�$�=�̶e�X�1�7�(��i}\�D�c]/1p�����<�q����%�g]���@v�8崦�j�7@�:��2���׎c�ݧ�קoiR1]y��';��
!|�KMt�O9Ʉ��d��O���)�$����I}k1�b+\%M����-*6��L�cU7��5���p<=�sMcG~�� g���S#�)Y�<��<<9��c1�#w��GL�#G ;s��[wU��uX����A>��w�<U�B�����b�pϢ3�15�p���;J�d\���<�f6�)�<�R2�҉,/A���K�sXK�[XxK���o�g��5���>�G��]�ה� -������Y.r�T�F<����������9����|F1^�8McXGs���֟�d'l�[j�LJV�ڻZ�6'a���{�I�=fG��sn�<c�7�e	c��wuc;����^�I�$�G���@E�Z+`�ET�0�NR�[2���c	(����8X�����x��	,G�f��/��ͧ�c�d|=�f}�ᬏ$y��T+�z�w�������
�.�1{,׫=�x 9-E�{�G�&��!C`��\n.�:�A��de�I#42�߄l���,X�zy'�Q*�a�du#J����w�<Q��~.V��UxP��Di�#�Q�͌�� ��?A�����޿�r�Y����!�D⛏V�� ��+a���؜�q��,�v[�8�ɦU�ה�,F����~���2�@�������^
1=��2=���#�7�|�.)ޞ�����7<4��S�d����=+�k_��k�o2}�}}ܛ���5o
��F������d��O�໱nL3��6�9���sՠAŞx��m��+؁��Ʃ�:t%V�w/����-��v�&�U��Z�W7d�\��q�ݬ�i�vi��tT���hD�j�G��]4��v���2Q���R��-�M����Al7X��G]���9�X&b쵤bM�iJ5pY��Id�:G�bݺ�Ӄ+����nVw��ʆ�5H�DĽ�W��Tv��n�m۬vꗰ	���YK�;���]d^����6q���;��Ǻ�h�2�=�AoS9�� ܦ46^���[(q+���^lq]��c��Q{StrH���@2�e��
�XJ�y�ן���/Oq����g��Q��懇��$�D֎���Ñ`�M|�iK�^��]B�	l||�w�'m�!��%bg�g�ςǩ�]�Ʉ��	��KP���pw0����3���NCѼ2Y�F�v�O4<�|�[
�ѵ
R��F��!�������;����8�k�ɁĴ+d���'�����k(g�ۮ���8�[/V��9�&�F���On��8�T�$�2�%���9^j�Q���a|��3�_i�K >
R<��oyt.
���c���`�|����1��2���G�{n|�tOP}��>�}���
��h��t�͹������G��p�3�A���6l�d��}Mf�]�k��{�7Dt�ԏs��cޟB0�#�?3$�^�1��k!��l�9�>,zG��vgrI�T��nZ�	UCFOk1����jH�JVb��#�Ɛ�;�|e���.ۖY����w�<������ïxg"�&��`s1�f<IIz�̾�����lV��uyPr�+��Uv�.��<|�6�h��~hdwY�ϙ���;L�F�� �.v�m�+�u��L�d�&�w��R�L��R�N5�7O�=��Κ0d���jO|R=c׏���eh��ؠ�R9]�� �q(lG}��-z׃�ݏ��{�3�m��:-��lv�k��\G�R�["xT�,C�U���u��F�D�	�_O�l�"�Օo+��W��q��"!�(w2��]a����t��m	HѰ�������u�����WP�&p[�z��s�w���U�J�j�Aַ�_���~=����8��ڧ�(l2�{�G��#��/H���s���Ԟ�ɸ���}n���n�����c>��%%��`)jv�ef�A�Gx���;�}>�Ry��jvC����j�ƾk�y������?	g��c���?Ci폁��4�7���R<��-��.
�����yB�|n|�p�������)Gx��(K�Ulǐ�-��U��,�ҍ( ��V3����3G,�Ċ�����K*��E� rP��'�wx౑�%�c�yW9�<�yٹ#i���Ө��\U0�Q\K-t4��c�{<�!��8�A�F��OF�
>��yP�#�b�DW�7�%���~_f|�a��rv�ZA�2�A�Z�mJ�;����(����f<��m��;V9b��e*d��m�߁�R?|�%�n���6*AjT��7��qDW�I���ҷT�s���m��v+;ө0�iemt
�fcy��Q��M���9������,#�B)G �xh��i��ϰCY�e)0iQItm:�V�����c�۔׮�]���I����`k�J4r�mr��DX�㿁m�a~���\�]�<�[�Z�H�-�E�x"-ot�;��
�^�[����8��SiT��D��R�!2*��mz�}�0i���,�>F�@��h��u��]tYK?q��R�C@8�a��Κ�9�Q�&�i��X	Y�e�����jmWhH>u|*��B�S�R���n������<���<�]��x.��j=�Lu�����K�������	�f��`9M6\[������O���zrX2�dTS|%�g�J�wq�G��.N~Ȱ���<����1h,E8���f���5����]��,��@�kʛ�kb�2�
H��6�)#bU�3�j:�FC�ۗ1Q�2����R���)	���#����k�p�d��K� �WG����C�9�,s��I��o��<�ò�C������n���H@�?8��e�d䪺��X	��.TC�]�cʻ��,đ���mA��9^�I��-ӽi4�_3���8�bǛJΖ���A��T7�o����G�O\oC�Qұ��#9N�SI�߮�SD{�F把��������Ƒ��M+����x{�T�o[���oA���x��MN��q�J��:;	c���Ec���.����� �v:J�x�X�`5�������ھq����+nE�zx�q-:Fm�L�-�z������gs��a����ʫ(�T�	�ä��a�e&��yW9�c�>c�:2{+����D'fx j�bp�s(&�B�
2_^$ib��s�Y{~��I;*xĚ)Z����m�:����۫m2q��0�[m]4b}�ۤk��\����^[���ݩe�t��$����޺�l�I�2�9v�t���-�f�+�|>x��m�ʩX#�:�E @�X\�{Ž.qĐu�%�}�z��[0�pu:9,X8w�*b�G7Y��;%�k��;���ln��ٺ��Y��=��P��<o!~(����`m���Z�M0���gO��.ʱ����
��#Ekð,�Z��B���nzٟ>,<��6e�ʹ����Tō���&݃�l�6�Ǡx�ZCP�d��{b�R梡�gݽՋ=�zUPjKH�!q%#}��s`��՗PI����ۦۚ,z��ך1��k��m�\]{��o�&eu��z�f̯���H;Z���1)'vy�;JHl8;�:�M+u<��Z8�4곯�U��{u��\
Z�z���X&�V�N�5͘��<��0`��λ�3k��L�`ڱ��CNJ��r^^���l<����э��DrpV��v^��ƽ���kmc��wS@�J�p��+���-;���I뇻��-y׏�i����jwh�h�Զ���1g�c���7�K&O�׼�ۨY����\q�-�&�u���k�M{�%6��D�O��2��J�zq���hMZ2g�{܌46��A#1i����A����=+�����'�*��y`��(��wS%a�;.8�9idT�4�ֲw�e��=,�&<h��m���㊄ٵ/N�q0�0�R�1s�v4�Ӵ���8�N�h�rGj�]%[<n��ZcD$�<ƐR"Ҧ���� N�t���M�]<i��M��Α7m�gs��X�궗v���"��N��n+$���Tw��o�A���}PMm80,�q��3}�(���KEhV��5�in��6y�,�k�r���OAH&�C�ɍ�Fɐ{W� l��O��M,�ײŤ�r�����n���D����PԽ�({��7w���������^�6�^��M�C0�vdq�;-lx��p���T,�Ce�\n�B ��h-�ހ��֔%��L.��ׁ(FL�b�nS
�o�]D,Tⅽ���V��&s�]>�xi�4Ī�u������)o�#�����q��-Ÿ�e#�Au�'_N^���橖Z0�R���� FI�z+;T��!ذgwd���-qB�.x�hY�	�G����vk5��;�거&3u�nv*�&�#�v�ݎ��/F�2ƣn�^f5� .�y�R哩�8ѹ�WTc]�ɮ{C�ej��4�F�>�Vc�5�t�1��P�1�5�ynP�tК��ۃ���;��d0�h��G��s����H��#�"��C�i�tE��'u`��k)X���\�)t�p�(� �<l�u�vU�s���;b�d�襗Mp�p�U.�5�x@�{v0��M�t[�V��^�6N��yq���{*��L�s2?nZ��dkp{#z��d٫K n�1HW,.L�8�ʶ�bˈ�n�h
!�i$�n^.s�,��A̅gᥚ\k<��ʹw����1�z�u�e#�U�Rbwosm|)#�@�qa��HX��	��i��ۚ� n'��L6�*����i	;6�CM���aB�Ir�XL;G���\hR��zr�_]9ɺT�4�b8��0ܜ����ѺfZ��jL��wm�U(g{ɏt#v�8����ā�T��R<��9�F�kܨ�n<-�(ri[�@6y�4q�B��{�Qȵ;�I�*�ءe�z-��}�~�;��c(�8kN��o�sjj�E��S������nOj�&�6:�,kP�[�8��/�W4Re�u[S�G-�h�c����K\���n�^��=~
��,�>P	�n�r \�R�}<M<�6U]�h�uc>K劻���Q�r�MY�0�������7,�'�^Ϸ�Um�dmMK(�r����E�R�Q<�޺a�8���v��={�KJl�\�t�����g�X�c^�6�͐X�u>���;��G���B�������(��A��U�Y���y�o��*��ug��4\k��/#K�����-΢�IΗ ;�6��'���ҋu.០k�-��7�O�Z�x�ܦ�I�=>��#gn�P&��7x������q�ٜ4MX�E�\�6�k Iw!��|�ǻ�����u�Â�3;�v�"M`��Fr�s��M�;¤�|+��XQ沒h�ę�X"w��:G�q߲�A��6�U��b��9v4�[`5�����s38X�'����SjZ��>&���ä5�6J���T���Ǜ��EB��i����],C�m\/���J��P%NYQH;5��w�����漦z��.�-�7P��~l�����liV��ffy�x�A�/�l�X�i�wh��s��u�����kr��0+�N�Bʵ�(]�`���7m3��=��S��'�s�Q���ޢa�φ&庥1�K�Hx͇�W���r��#:)g}X�{u/��C�Wld+vP���E���$�QީLex.-��O��3����En�n1^�t��e����z�*(�>NZ:�E낡�E��:��y�ݾ���:g�j�rU)$��K�F��ݷ���&������YL�֭t=�shP���i��p�'#��;lV;e���l�_1��4�o|>L���[�Q�{�ѥ��{�w�l����/�k_�Yx� ��Z��匝�Ȅ�,���`�Yu�_���J������kY�3R�j,��S��%�dEѸ�θYY���N�y�y��-��y�_�<\
Cz��b�k�ͺ���[rk]���J���mAٯ=&�sВ� x���wT���1�d_0:�����;��a�e�J>{5CF����9��u'�w�nnza��P�ʕA�v{�����R�Ƨ^O^W���k�����]��/���E�����=��!}��~;I9#~������V9fD8���/%1���p��7�z���m5�%;NI���,�����վx�^�Ǿo���Vo��>�ݘ;�«l��J��c��pٵ,�W@�5��j���#W�����m���P#.�\��-a�.���<:�w����	�kXT@ˋ㟕M���A� l=y����u��90X��v�!���YZ�6�i������ǅ�Ӻq�>�؅�l����)�=QR,����c�j�(��M�ဳt�А@��n���}�{��A1)�ޕ�K�4�u[q���L8���<���A�U�
���+�k�k'x�M�5v3���c�K�M��z�ݮM�Zu��O��%�YY;F9�g؋(H5�W��nj|�񶆏Zce�û�+t����*Dт��]����}�7�wP�g��':D���8��W'�cǋ�n�J�jm�ʹ�8 eƈ�����j����H�/p�eA�gm{Ƞ���M�y�p��m�=q5�871�϶#a�Lj��fCe��yu�Լ[��ڠ��p�p6�������=x�K��e��î-g�@r��=$f!��%����qZ�ٌI�.^��Z�{����%q�$��2fs5���&:�n��{͞gް��_���v���aX<;�ҝhs��qDA���<p�&����������R~]��պ\R�-%l��+e׺*<��Ý�Qx��ڪԃ�B��:כ6����G6�:���fg���6l�;�Dc)ɓl�;խT��ƀ�o�2����%u?ќ}��˕9T�"�Pnˋ1\N�dq�U�#6��b�A7.�2|�ũI�q����:H��y��<c�ͣ:"-�T����ƨ��n
��eo���pZ�3���-+�)�tj��7��}�T�>)j1�ꝥ�6޻@���v������tg�S�[*$�eadD�O�5#h]S�xxq�p�CHI:rQw&,���P��Y�e�JR�m�)�l�;[ m�2XMQk';�Գ�v��;���b��'$of��[�E��,nr�k���5��,
�`��_1��d�l�zZޛ��4�#lzg)8���,��9��!D�v�oI���Mv��Ӂ�t[���>�U�U6�5���{�0�'����):M�ޝ׆f�m%�Ɇ���$mJ�p��,�I��l��dW���>j3�����f��ӆ�zQ���=���<kI�����E���|�76�6�N݋��NVݲ,�y��Kg]���}�<��Y�&���6K��s��g������e�;UM�h��E���H�m�{�y֓�/5������H�
Z�"�.�gb2�6�K[���>�p6u)�;
}7�H�c b����Ԧg�G����^���15�L��f�e1r���w<�S[AT��f��80�����H��-�:�����Z=�s�4���9�Q*b�x`a���|���}����٧̷Ȗ����q�����fL�B�r����z,�2)�b�l���;,R���>��(�~ith"Sj|��(D�9�S�d�[��D����t1�����5��g�N��a�d@42�Ϩ�����JY@�r��[A�Gb�r[/CWK^Ir�V�kt;����z�������nD���^���ո��Zzy��z��A4Fkz�;���=q�����#
�nn�|�Gv�:�b�F�2�Jd�p�oO@Zʽ����[7Rujj�8[E�S�����p<������:��e��ǕCnͫ��d�v�s�/n�`P�>��mǬ��`X�(wT[!�¯hu�v�]����vy��[�E��#���;v��0	��vh�FՊ�G����S��������H�kTY\����7+u�H�����>u� Ҟ�Y<1�u�$�t�|� �lč��KX�3���sv1Fp�� �l����фE1xHXH����< �%�JR���>3Z�)+˗TM_������3D9��>;���Q,���y���$��shd(�8�E�ctZbca�9���w"a�cJ4���r�����:=���r#��Q�*�Q����ΡEox0�&a�nW��j�R}�L�u
��.־�k1b����>�[lqϳ�5��<�Xﹸz7kUX�T*!9IvyT*�"H��X���9���_��C�Qʇ{�`�ņ#��Ur~S�ah�2<wT�w�y���2�;��Gj�M��	�V̜;39!h��S-r˯pǟ������-q<�U0�m����q�g����X�U��)�h2�D�����ojS�c@8i�p�D�1}5��ݨa��]Ŀ����:B���9�e���M�{:�'w�t��Ñ����V��d��{Ms�Ɂ�^a�b�=S63��1�K�q,�Ͻ��d����K.�q�P���QKnA��md��;t�֩�c�����qK�Ipo��3�e]�,�g�.�@�n'����x�C �΅;\�^O
� �|Φ�6Y�1&2�b��:��t�b�j����[r׺^��p��U���olt���N�m�՚��H����Ν�����|�|0Oj.͞.J砊��[ j�:8�3�V ��+���m��Z�W��uݒ������ur
��8=Nޢû�0E�GDJ�Ka]n���{��'��\��.��j@�6>t��2�3!5,'���G2�OD�̋�!�:Ĵ����\u�xU���L�eX#H�N+m�8d�X,�(ⶀ2�]��$r�ϟ>���q�P ����#L2�������;+^U��J�=�B��,�~�:�R�x���b6֜ΎE��3 ]�Q�9SvE#�ۯtY~�b/J�圵�{5�Z��Ɩ��,"qut�w1`u�Ri����R�[q�ȘmF�:����:�����������Tv���ȄP�5�稨(����b�@.uچH�\�,��'qQ�xLȼ��Ï2��y�yw#mW�k��7'vcm�z)�`�x�[l�Mf��|�
�_���\M!R[��Ҏa!J�j�)���^P33lGC�͇l��8�7R�z�:�����L�5�:\���ɝ��@i�v�8��K=�m�y�y^@�%���ˬ~=��~:e�p�}ܱ�8اn�,�lt���"�݃���Z[�F����r��n}�&�i=j#���A�'d���#'&c1�CI�5�g�3��f�Nlv�C_��x����]]F��u, U0�l�ny�l��I\mV9�$���V���䫘���T��\{D�1q��`A<W'ז�(���2���J���p�`�{���������C�T��lD;3��h�
]��Ɲ���md#K�_ �#_�d���CgOH��|.��ww���#�$;��8^݂���qݸؘ0�Gý�%�!�V����ա�kzh�z�Z��@���}�� ��HN����A������ظՒ��t����{X���M�wl���Sz��a�j��n|���1f�#�8f��/�5&�v��4�-�2����@�k!tYP��Xhmã��|�쳡gLDx����JfS���l���cL�w�",bH��+L����s�ң̚��;�xYx)��$5Ƕ��H(��ٕ���](w �"��3���N#R�����XZ��\�"��n ���DY��a��&f|<N�:��g�x�#18���Ⱦ�9s���?A��ӈ�
;j����ɪ׾6�>����lb�6<��.�6ƕV�mT���n�z�"��*W��G>$P��ё�MTڅ<���<,�朦xs���!�쑧Gp��m�YP��^y��|�����;���������E�s��1�|b����U�ޑK:�x�"qsY�ms|&Is�|�%5�"қx�w��Z!�7���<7�
��f��n�dc���kˎ�Hm�E�M��W���s�9���u�*��6��ڙC� ����&�pP:�.�R8�*Q�O3�M˵H8yũI����M��}����Uj���\R��Y`��\�{���|�2�>I��@�p��횕,Wb���v���1�՟ <���l�Lrg���ԅ[��N�3g[_vV�����g��(V([j�Tږ�]-"YW��7y�x��i]�\�Ɇ��x��CF�\t%���[�%��t�ˡx��x{�� A؃:ㇻXI�P<G3��Gj�	�]� �+���f �dB)�p��OZ�x���n΢y`�a�� n�M�8�j���J�予h��ơ	�;X���p�Pױ:��W�t�Ak <;�QF�1y4cq`�N�YH:���\P�5����)���T�}4�܃�wJa��\o�����	����.<n�ƥV�:��3A>�EV�g]�Œ�&�!\՗U����gz�f��=��p͝��ió۩eҧ�F�\b�:�ٗ��&�H@e�.e����ݽ��`��Mm�������]�4���s�M/I���3�e@rwE�<W�D����Z؃�㈰ ��q���l�+"�R�kjນ��y�;�l����㹛m�K4!Ǌ�~�$�9g.0��9 {�d[PWu�9�xծ�Ec� ��z]�/KNǟ�oSj���?"��QT���|�fe<e��!�e)L�����"���7<������C�7M��ƙ��{ܘb�4G���٨c2Z�w6<j��e��ޤw�9�5ֹ¥���ӄV�BZR"R@�k�6�~H��r}������(��X�> �i8 �"��c<P��۹*�?FC˱�K��<T�͸B ]F]{��\��x<d��f<9�Y7�.(�d��Z�v�u����=u�b�4ufށ*�;��������n�/���0[we2l��g��q�R�/]���溛���u$���[^2�bk���<�X'x����&�;q���+
o:��<��Wn�ϲ2�^ZF�o"�,�����a)�_�5��;3�	�5*���P�&]�c�يQ�X^���T�'+?�E$鼏�h{��wМ�.	�M�-"C�����>����܉b��������m=��l�^�)��wq���F>򎝗�(�݈��L�3E�Ʋ1	���,��|-���u�R-�u
=R��,��]���(�\a���VR8ܡ�9�v����n�3ۜi۔��S���Ba��m��k�va%k5��2v6#�H����s�v���'3ꧭ�ɍ��m�˭E�pF��j:57V�2w��Ξ�^��wR&�8�SX3�mip�6��s���z�9p�[v����[0&�h.dr�]KL{r<v�Ǟ�=C�m<�p��q"rp��mqSn����$�ó.���{�`�bm��S:jVČ��XI+hO6��xxi7�j����b� ��/# �m|��>����~H+�-*��Qg/#�A�d�i%e"���F������_�!^�i�q'{��g�N넞��1}_MN֌�p�����X��H\���pdH,�5 0|!�˻�p�w���p/�_�0�y �C�J�EVf�X����}�u� Lh�@y����S�D�~n�����"�� 4�!ϙ�8���ؽ�����M��I+N�VR��m�H䚠]�yD�؏*8&����6�ḍ��ɨ�^|����׵�8��f�*)pՌ���~D�[k������G�j�.�2�3���x�*:܊�O>�8�(�����������?��Kj�V����؂�	�0����_|J��im��5;�!�@����v�j|�^���79v��m�8��n-)�����t� �#�������&����^�x�������,������#v�k;{�<q�=�8�y����i��Pӭ��	Ӑ�A�=]dv@�Ok{���.��v1�%�u��8���"J��"v�F�K�&yC2��M+�����yT�Q�Gy��qR�{���fy �n�!�c�w-��,���%��R������@t�����5�y9��bQ�H��ݓ���,/6���&�6ƫkh�TF������*W�K>w649�4ޒ4	����;�m'k|���W{f`��>�S�m7R�j.��p��1��Dv7z������z����-�Vm����9N1�Gv��w2�%�v����H���
��Ds����(n����;���@�O9�2�Pu�xC���˟x�y�l�K>�ף�I V�X&[m�]�Z��G�=�	�q�3�򝎿!l=.�5�����++T�^�n$i�U�Ey�y��P��4w�h�U���zm�{/�^�wJ
X�fN�t��I��0�&Y�̐�[U 눦��><�әU�H�k|�th���|�kl��v;F�ֲ4�c>�6@�>Xާ��8�y��֪���Wkqщ��F��DI�{�Ҹ���v�sǜϼwU�w=��+Ð�ܕ�����Yu͑[�/DT���>߀૶\��άd�8������a��X+T
N哼�/q�4WU��Y�� KrỮ�6@��7��|i�E��A�h�ͳ�̣��v��9�X}�x4��ݻ-��ӌ��&��ج�)Bw,��E��{#ڴ�p`Sk�^����v,���͡����7*@WbʚX]L�x�=s��9wzM3v3b�\���u�5~)Jg�^<{�q�%،�ƀ�j#\:��3[�\4�5]�F��-?|}�/k�'�����-T��,�Bu(t����6=�[���b=�lK�bw�s-a�î��h^�@�7��P��e��"�N��=��8����K�ϡ&�YZ)*�(׬�؜�`k#z�x��{��v��ci������(}�'�o"�3�ƫ���!5Xf��2����Ì0Z�7`�^�>��zq��xf-�����kӊ��oQ��m�'�3F@�k����_]*{ޡp!�tv��E�����������/�}۾�֥z�̉��X:H�f;FQ�S��d��������/�^�6=��uN��0�Z�,�e�Y�6�9���'<e��p��[����21�Rҗ.��_��h��6���¶�/�5~Z�ơ�b�G�;fv*���}�;꫍V��<%�Ù�����d�V�����*�Q� �d,�3��l�k�7Ǟ	�}�C��)��5�� x���{eO,'D6��8@Ϩ8���@d���Ԍ��
;}�k��'�u�צ�S^�c+�vF=4z����G�p%ۍ�³sMm�(�B�ۉ�	%�����$�w��ǥ۶�[8���
##��n.!�ϩR�֥+�C^f�>'��jY�8��n����)f}#�˹��1�x�.+U�V?PI�k��və�!���\��̂�����4:��˽�8�l�_��HUl� E��!k ��֡Dn ��cd9�R��Q���Ƒ�%QFw�x�ɥq�h�m��@#uY�,S�tlj�7a���F`��>ߟ���aHa#&ٷmE�lC�%B�\��]�͡��-��st������k�����!�`�%�CSGm[B�0jYȤv�}ƫ��J�k����L��fޓ*�;���M.��v1cխi�2۫�������P<�s�8%��e-	��/<�xMm�}�?�8S=k�d�~���C7ۭ�f0eI�[����������q*<�P�ܠ [��b3�M���5�m$�Ե����(��E
����=l�|s��:�CNdy�{1�"bʆ5U ��~([∂2f�d�Dʼµ7t��1(w�����>��sq`��;��.,n�%���Y�V��(����yK�;���ɺy̹�̀��F�V�^��.Ό���r���b��!71���;��xw%Q�n�'����x	+�ܒ 7TTCn��r[��{�G��[���<������<��qR��Q޵ŞH�7S�Ե�%)��r=�ٵ�[��ɂy��Y@S�^YA�&,�`�=t�Q�!ㇵ٫��!���޹����K�ۂ8����==-���ͻ\�l@/kߋ���)�{�^�d���T��yQ�ɢ�����&���5]�F�4�v�GsdX �+���9��i�M64��W����8��Z�j&�d�<�\���Mt��ir�%�"r>T�^�M3�|�9��U{����.�
��0�@yA��ީJ�;��N˄�����c"�
��(Ymz�m����M��xu�L�by�����W�Dʚiv��v�d�8��ׇ!Fa��c|1Q����)f,�kǈ�y�;���[+�RX܊�%(��q{����L�f׃q�E�yĪ/��߀<EZ��� �Dq���Yuu�
���E�h��U�2��8��n;yKX�//)X�Ѧ�n-,��Ύ�(�~6��W��%��l#:�HsC�uY�s\"��A�r�	M�\� �՞�_�s}�|A#�r$�I$�P@(��QP@>�5�G���m3��&"Xq��Uܭva�%��%���� -�� "'�7��TA�Ie �UD͊A$dA$$�2��¥�	+". �@IY�I$� �G,�Kh(b*%DVE(� ��� ��AB��(�b
@[PB� Ej ���&����&Y�h%���$'(  $��
� ����O����m2�4ϛowI��nm?�r�8�����jbvC��းr!�7��=_��~ڼ�oXG1܅�G0y�wt��uu<{C��p��s��`d1�����_�����{@@5A �|����G��������`{F�P��|=�)����d��T'���H��C��Z{�=�y��؍P��C�{aE��.�J��c,�@=O7@L4s���-@~����v�dEX�Q!H�@R$!�	IH�Q"�#H A*�Q �Q"�D�@(�B*��B+ H�"�H�@��
0"���"�@�,
��@�0 $����$`� 0  �"+""�
*�(� "+*0 �
� ,"@���"��"� 0 ���@�@����"���@��@���0"�@�*����@�$�@��"$�"��bF$	@�Dt` �яB�	k-;�l�fw����'��ϵJC�����������Q�N�2�j<F���|#���F���#�����h"*����|�q�������w�d \:����m����!a:55�Wo�p�v�����ل��ɷ�3�}�I�w"��o�'�������u믮m��:�ה E �X�EA ��z1}Fl�6��`�j�v@<����x����8� "�!�C2������aO�&�>���3��l�(�J�a�L�p.\(2/h9�P@%��fC�z{�'U�P@:���A�9��D*/�~�p�/4�`�8�_*u�S����|����E���K
��MD|F���܊��8@:�?Ӈ-�O_��7NC��#� �x4��)�6w��;̈�q�����i�+���1r�jm���� ���U<�3�ڞwa쁡�@�s /�1g���r ��{�����Ȁ��h|���/$�<��EP@:�-Ґ=�sK��<s���� ����_(0������w$S�	��