BZh91AY&SY@1[�_�py����������a%� @       @      
 g=*%

��UP�@ (�%U(PE(�z�P�TQ@*�

(�� @    ��@���
������c�ݜ�^�{���Gѽ�_O{�� �ѻ�B@�P��E# ފ89���2@oc�oUG ӟ`yl���ڂy
�G} 
��C��{�"�C!�I����UæX��d5����@(tJI@��h����x$�c����H���H�0:�)Ep������CF�^@p�\� ���=^ۃO{GQT��Ug ^��:pttt4�	�l}�Z��g��B�$ �+GCL�]�;8t}�zh�X���m��@T�*;���{Αű���v��0h�݂A֨�E#y@�����	�A�N�0����A�OKc���P(�g{� �n4hd�e�v����t1��9���� �@ �� P  �  T�2T�P�@� � CFO�Ĕ��р F 0 Oɪ���R   @   ��JH��OSC#L����&`�OT�i5P �� ���  $"4TMi1�T�S�R~T�6�4�@{�16��S�}G����ۿ�_u�O��A ��j�� ���P �� ������/���?���zH�� F���UJS���� z�M�8%1E ܨ����a������؈(���_���]g��K�t�]�w���M�~�+U�سf��&�A������,���=��>�R3��J�K�U�)����]�}�U�Ge�����8�pP��پ^ۛ�Sק���ڮ�s��A����Ξߴ��T�6�*��e�-]��T3����Ò��
?�L?|�
?����W�|_��B��,K��j�ը+*K�)
+F�>��f���হJ��2�.Ĺѹ;����s�$5mh}����X���i����͈7�IU�� ���1.8b��P87��2�i��:{�S��6�P�Aa������tX�=gD�p��۱��m��?[�Z��1��i���FI��5�]����솲T�Sn8y���]��Ȱ�3t0�'�K�3&ûhP#���T��&��x�.܋�f�(^�#�aܗ%Z��(ŶrC�fl0����>�n�n�N����6�9��\ذ�� 0@��wH#��L��rX�M���3 S�R,�s��R���������j��D��o%:��a��3V����075��n�]���F&@*�x���*0�Y��}��
b����K �u��"u뷰���wI��U�6kۚ`�F����ذ�1؜"�@Q��p��������U�e8�ަ�:3�k:zGEɂ�k����n�CH۝#���,�aq�<����Gxh��4�Ҥ��j�dx���⯅tkE��{z�l����rd�Aw��q8�i3`��7�c�q�	䜊�F��0ؾzW�F�ת�Mz*r��,�
n����0sF�^���#�����gM3r�A�N2�ĺk�ƥ�x�]�֚�;�X{ �7�o^G���S�����s"S-M��ڳN��^K�b�+0!q�94,;��m��O�Lm]Q�H�*hrG{B��wۨ��v1�B����%�m����.1�E����#�T���.]�,s������M�D�uX�Gܳt�oeY���J/7K� c�s�t�N�kmốh�Ǘ'�3�Y��7;{�Ca���٩����(����4wr\ڡk5�U37�1qi���m��<LջǶ�f��pWL	q����/���l����է��2��./�tmю���C�a�%n�%����m�y��9������d��K�����eiǗ9��X�^�Xl�����V�;�{��O}��m�(ŀ�S�A�GЎ���6�ʐ5��a�����G���;zC�>Q�F٬�ݔ�W��U������Ԏ���;���mN	Ō�l�N�Xn�E<�k�h��T��D������ӯm�5�zu3yc��y�����u�a��
�(�e����c��`��ɠ�P9��$�ݛb��mh��k��=-��K[��ley�ͫGe��\�U�D.kr��xD�����YT�������t�Cs��3t l9z6��꣌z�Nǀ���!tҧ��5�āi���yХAn��3D������(ƺ��oǫ�Pa���`�9*9{G{Y/g-���U�1~�@5 ��~�lR�hM^�J�x�\U�hѫz͘c+�T��+{��#Q晃����:w]Τ�Dّ���ѹ:ՔnI�T�Ҧ�&�>�vѷ�E�$�0��F�ޛ���LC�% ��j�i�b��:-�T�;��M�jޘQ
���L׉���{I�Kf��N{4n�ɦ;k���G��]�ݛX�������bkp�t��9���/P��G=Ӏs�Yđ����CB�c�N��@��ڹ��+ѿ�fh�6��a�����M7zn��h���L0��k�Rjv���rfm�/o�D=Mf[�:҇N�(λd�����1�����=��M
��)��8`�1m�b6��wh��p2�:�N^�)��z7�<%�k�s/; ɲ�-�c�f�E�o���_.ԮuZ�m���b�%��~]]x&�s��FN��̋O���o���ym��Q�7���Ohs{�p����C���"Ɉu�еb[���f�N���T�+*x�-K�[���7���Vu����3�6'���"V0񐐰��d�B�D��7]%�������x��Kn�e��^9�`>7�K��gO��O9�>y�,˽�oJ�WB}b"�X����A���\G�7Ε�g�����4�C>���!���z��9q2�l��.:PPtѷY�t,b�&�B�&#�]oB��R*ҥw�;{p�����O�f�9�p�w�;zl�X ���x+K����Qb=TFi�6,��H\�\<��`)X���[$��S.�jhbހ��1�}�a�=#��3�n�\�L�f>2E9���1�$�m����I�A\�.Ϋ��ڻ凰O?��
��tX����vԸ��ur�!�I]�^���K^s�����N�&��Bܐ���E�zK�Wc2-�d�%L�IChƻ�{��읇ww��ge��i�I!���Q�Y����9�hꖅ^����`���h���n� <�_�촗�7z�{��7nYy��թ�i�L<�������:���C���'wI#WkWf�q��Q�av�Z�{��2�����LN�C���":K�ׄR�woS�W�b7
t�E6S 8u��8֌��9�Y�l_J�]�-ڧ7����wL�\�v��5212Ҷ39;�&��h�gL�J�C�x���Np����z��ph��p�C�nt�qB���곋�,�`w=���Y��`Kz�x�=��ùǉ�1tH�U�ԫ;����*����T���������-;��p�&�P��|��ag&v����7����%F4n��8橌cف����FA��+(�U��!Fd�*,�7�� pf-L>�ޜQ�5��Z�a�;:�NO�c�wN�@,�Q�oC_5�u:����WL�3���d�v��*��ggU6\����6��p��t��Y{�����y�	ڸ�+2�;�Iǧ>�,�G~-�E�pe�c����u��AC�J��u ,$0һO��/�V�^8阌�p��\F���\��x��V�Sy�]��5Vq�x�rma6��� A��AF`�h�� �Vk&��Hqwu��1�W_=�a�	<�̢vn�x٣~7/L�œ.�޷WD�6�s����iY�����Թ�8	Ǘ�r��*�]�&Φk�3F�Ku�X�NT��Cw���}���0�>ۆ�Yk�;�ί�ɿI�1��wg�&�H8LS9͚�L@�<���L��\V,("p��&�"O�oo/��
M,�n��w�>➽��/f�j76�#�
B���ŭ�B�bߞ��	����&�\D�����YA�BA��<�c�ـc��\�Y��$����D�яF�MS꺹Ӳ���s�+�i�J��'Ln��MbY{� �J�̈��K�W�A����������v��;�b����ծ<���&��� ҂�ni��f*9����/(�QF��lZ�F$k3�0���E��\C�&��v���} X��ꦨ��&.�.v��:^E !�8$s:Q�%�uQg�sMכ*`�S�k-f��{�<p��f�h�;���~=��q��r㷈��������#��uŔ�oZ}�f��4'�3N��ur[��;0�1�@Z��0w	B#z�Z�{�\Rh�Hs��ώ^�'63P�~�>����
�������+����(����p��77����ﰨꟛ����0����&��ʓ�ˆTo0nvو��M���v�ٮ�|h��{8��g���p˱+Z3%x��b�ټ0F�k���_��p������4�My�ڌ�Îu�mp&��wGHgp��c�\�XKu�F�x��Aёͱ��QM۞��������-]�!�gV�el����&�6+�3v,��[E{W\ṕ�e�x��lZ2��<�F�7v�4%�۬#�A�ugb���U�J���AeaJ	�]�Utw+6ف{T�M�Ȩ��:�,h�ˋ�e��8?�n���mڰ�Y�ϕ���Uv킽�}=�|9���<vNٹ^���k��6�ū��H���z�t+b=��p��ۭ��v���t:s��v�<蚺�sm[�1��K�Gq�%�c:��e�u�.%cB��9��ejۊ܆Ri]taL͂$o,�ҍVۛ��w.ֽ�6�%m`s��ٮkn��ѭ�[���T�,eц�/-35U�(喭�k�]����#��:���'�xE���T�WbgZ�;m��8��Y����nѻv,cM�ˊa�\��6E�$ffכsI�]f�`�b�6��F��6�ڌnƟW��Gh��S��՝c�Eܚ�x-�#��,��i�s����ɗmu�b�A�س��3:����c]KRf�l�!�1�$ֲ݉����
�\k�n7?/�����45�0�Cb�i]���RZ〈1��w%T�F�HD��kK�ǀ5�X{����H�^���Rk�����Z���N��Q�'G(�~w����}x��4܇-I�4�4��c�\CPp���(阍#��]BS\+6k�x*�dn�7[hG#v�Se���+�.���ZƘ��·Q�<L�\9�k���i��������2��JǷ��9ѣ��^.:��)����`�v�33e�u�H�3��n�+r�{���|0�ܗN4%�8}v+��R�u=���^��k��ĥ4n%0C7���m�u�p�⋲��;�;b�&��v�����@�68����R���\�,��]4�t��S3Y�6��c.xX�]k�gY�1�!����E��i+]8���m�1�y��X�Eb�a�����w�[�v1�s�^�e^�xy��;�@D�9!�G1�v�[h^9�q\H��t;	`�š����{&ۤ�M�֎���6�X�O��Z�ɜù�U0]{��N:.ch
e��Rl��y�#�f�����c��\�I�//jnN�-�휊^j��|qEm�e<���&�j:���Y[u�+�t���󈪺6D�l\3՗2ؔZ�k@��[f�[�fÝ�z�K:)7q�x�t�t핂v�1��sݻh9���Μr&���V��L�6s�=lK�&����m���\f��F��̧!�۠�I�0�o6�uӶ��n.��'E m�����#͉;M�[X�u��u�I��^�5��#v,���HT�C�ێ�	�n�t�a.�n��jc�Kᫍ��p�b6�˕�V�q!lX5烥�1�˯;��Y�]��.���\���Av�᷋�p뒴��nָ�cn:�m�,�q&ΔO4!<;��rh��{�ml�&&j�i�-RY�a.���j&K2-�R[��*��ٸ�����3O�`�Ρźm8�����I��֬;�櫫�a����Gi��ړ5�Ef�i��L��w�ъ;^j^�����]�l���;��iyr(d��\�:�b�0��jbkf�f�1��.��%Z����#ɕ0]�v�z�U�et���HC1��5���ح<i��bC���:�1Y/O^�ڍ5�[������A��mq<��ŝxw^<=3Π0v�����/b�� ��m���Zx��L�q�w)�װ:1Ln�V�e��Y.dL���Ɔ���s�GFL�C�E��ޢ;�o	#��u�������g[cD��%���=vt7��d ���x�F�m�,n����:�b���s%���U�h�V�z�F <�'q��&��Gvֳf�2ܑV�������P)����6�km@Q��谲���Ǉ�=s�+U�g��;2�Ob��<i�uqy�K�� �ݭ�J��+�V��9�������O�m`�=��Ό@m��T6�l#��T"��\�s����q�\xs0��H\������U�D�;����bd�;�jf��;>7K��ϋ[�׀���:i)�4�f�$l�7Gj����9�z��nJMs�ʙ�2�s�c89��I%fn9�qM+s��w]���G^���d�)�K��eUFd6����M�k������9����SEn݉W>�.(����#���u���6y0�WGO��Nv;n
��>@�:	}�N:�׍�kE�a�����hj����q�f[q�]Tj�[z��8z���6z�cQ��Sr�͎ٓ����]�qjV)4�x�g�9z-ק�GY��GN\ܴH��:*�,Ҧk�η`�A]�M|N���T��@��;P���ITN.k��Kv�k`�]���ΉR*Y�X�趬��ͱ��̾�wv��ml]yF�WL犉��i���<wl���6B�cm���j���Ѣ��֍�5v��4,��<���Xm�dh5j�n �n�ۍ������l-��[���L:�\�=v����i�,����̪�W�92H�`(��l�����UބC�7�?`_�~�>?����ߩM���e/�6c3M
pnzڲ �_u�� |��k,޹�sbsm=����H=ұ�1#e%rv&(N���¼��`���	���I�7D��M�|�rΐ?:/���~�p���ׁ3���'��A<��N�I���;놂�vA�y`��q�Y���3�0oTЀ4��j���Q&n�㳢����'���-��M����K�Z����Is�,����w'��n�LN��	������"������<���k�ni���������Ds�W��/'Hc�>ӽ�k~�@|������d݀=E�x��
��|q݌���a��f2a��'�e�M��+0�ظ�.�[�'��}Z�&��0������e���]����FH�=�P����Ky{�K���8g_��@���{���K����T��r�>^h�C`[�������lټ!WtƖ�5���[7��}��f����:���Og�t��w����ŭ�Ź��X���Z�E2NX@�,�����d��T,��x�6K��"�w��{xm�#'y�.�`��m����wþ�:�\�����h�	���!\i�����=��3^:{*F9Gp.��n����<�O��So���f{l����V{����d����k���wė�w��cW�a#�k�!|���(w��w�	�w���e��)h��^����`�
�b˸�"��uV����^YÅ�	��fW3����h�qϻ�~�.GQ��t��{ϓ���g/IW�n�]�s��=��kT+4w'Z��^��"a�����������s�3��o��+��r	{�xG�2�z;b��W���C��1�Iљ��t1y�z��#�Ó���o\ycȱ��/w\�rd̍AZ�e�[i=7�ٽ���^wF�iL���޾�G��]ΔXDZ��1���w�s�	,H��M��3��[�~�/6����g0c�6�nmn��bw,�59�N��؍�S��f�3z��7z�Ƿ��圲
������Ges�z��Y��y%v�ξdN�R�xhb�:���������Y�)T�D�lL��0���X���&�o|���0�}���p��]}f�E�0�G���E7N��vS{���]~��#���P�����o��V9��/sxN�ŏ+���.q`=����L�܆)	�t�f��������x��m�N���͏Ӊ���2}��;w���. kCI����Wu���>3�{����g��E�)?N^˰D-�T	�6pa�M���Ի�,��E.�k8����5���:�v\��gOz�?#پ�}����`��Y�x����tF1���g)��5͐��o{suމ=�Kc�U��g2`�/nV�}��pe����?N��Aݸ9���%6�ˈ͚�����9&��M�����i��T��U������H̔�ތt^�S�F��{�TJ��e�|Wxy�)y���s��9:��^88b#�����b��������:�z:��+[�^"�=}���x�:6��.������qz	#�9ؠ+�ۇ�v��z͙�F���S@jMc�Y,�F�gOo���4��{� �{`�����m�-������N������B����<�2{�j��s���Ux���:��!�9�D�7L�3}wt=zK��<�#��#�<��V��p=��oe�=/2e#x�'�r�{����B�����>������T3^XQ�Q�&�KH�C�ژ���
l{�,c7~����ú�Z����VqRy-}�6���j���<`���DtE�8{�wl����G��
=�A�׭^ޝ���f-n��f��]a&-}�5§��e�t,�����9�槕����eas����7�t�̸Ꝅ��������&��1���[����OW���2T���o����H㺛��;�!f�4h)��-Ƽ9[�,9�snZ�n@����X�^�Ps�oG�x�~�~üj	��0՛����7\�h�^��yBrl��{c��K�kx�g>��{��8���	��������E�ȧ�[X0rY�{����J`F�`�#�C����ۀ��/��q��٨A���^���9��#�����u��D�4I�cI�n���q��Ek6cB�8�V��%�ֺ�eHn��L�z=Wزq��f�@�ؓ�ڱ�+I�I:�y���j��[<��ػ�4WU�⢙�J��IVm��S����|!�𙷹?yz+v����vQ��U��8���U.{��Oc{�;�;�o�qܚA��?O0��G������{Zʻ���{g��d��w�j��-m�sv�ZV>߯�y�Z�1����ѝj�^������X�K���}�}z�����w��w��O��~���< �5q��)#w�d��6^�Vn����0f��H\N�|0dn=C�~>};'{<_x���>��	z���HaT��N5���`�'��{u��=��,�������]�M�}�[�Û��}}&�:M({Q���z�+u��gHZZ�5c�(�No������V=Nۗ�u��]86A<5���l�|�i�X�ذb��|Lٛ��J8}�1���{M����Rˢo�P�C��|���ҡ��R���l��}6w�)�W.�~�<�.O�oōU��=�ӯ�t��ʎW|�<�ĉ��j���;Ӧ<��{�Fsi��G)U�?!���ø�_<S(�m{�t��;��	Ҹ��HY.W�uY�wEA{6���.>ӯ��Ns��gt6Χ���7̈�kY�%.��ێw����b��h�3gx��
0Y�3PC�o�����V{ޣv��
���2B�S��K��&=��z�M��C�7p�7#��M�or���yzw�>�i&�r���3��"6�Ƹ�y�y���}��L�~�Y�(�Y��g���ЉW/,����f
��cp6��ɷW��×�ǣ�6t�T|��q?o���n{i����Vj�uh�\>]{�η��+-��f����!�{=G"�3w.v;�,�qn�Y�� ��P��B�f��g��Ճ
X��,��j�r����丼\��r���y�c�����:��z�E�V$�x������T��c���P�
�	:%��c=6�;���s�Ղ�K��o�]Ҭ��N�X��˼6� ��tC��y��2��FptO{=���K¶�H�_!�u���^>��v�|T��j��ŝ"g�ｇ)z�^ߔٝG���=�
�Y�\cq�o5��%���w`���`vɗ[�}o��n^{��g�޺��$��|��	ѳ=_��O�8隣z��-ܦ�<��B2P��X�޼[Ӱ�t�/��R�x���4L�3�q��]�ԺE�䙦��cވ�.Y}Ӗ;ɟ#��:Ʀ�4��t�f���>��dɣ8x]:��w��4(��u
�`��=��E<�MT=����4��{�(��	��	}����Py�_L�U�垊̜��.x�\�1��2����K|�rї{|6m�AB�W��I����Goy,��=~�0���f���u�E��ݗ�$ɸǷ�'����{�V֟�y���[�V�ӕ3=o���m�7������j�����s��s�h��Z�����;�C��>�}����Uy�T&��ɽ�1����yд{ُ%Ǿd.>��sF�ՑU�OW	�7�6���u_q���6��q}�g�.�m��W���a�ȿ����`S��| "�W���������(x�Ta?������;��,�H�y�w��;�K��42��e�9�;s/[�۫�l�ŵon��cb��əa��H1���f.YKp�hQ��1���#��s�"�E�3cj�8=r���;�q:^K��|�ٹ��\�Gb�r��]Xy������1��l���w7	sOf�{S���6�ٵR4�q̬Ǝ*�͎����ڧ�.�����1���e��]��������gg6�Kͤ�u�r��l�<��/XGG<�ωn��.��S�kZiv�Ux;pWknm�.����th�y;���;K��5�Y�4#@(3F �ȉ�I�����ص�f�Ѣ�hI�]�CQ3/`�J:[Z����.h�.�Ny�7v�;�k��;�K�_k��_��V��
r�&�ۈ3mΖ��2Z�	m`X�1ְu�D�RP��!��%�9����n�SS���1���:�e���m��QT`m��.���1��y���\T 쌵���736;f�Z�ܜ{Km�rE���qn���u��q���I���dJ�5A���Bһp��m6��-���j����__�;�=r���~ζ�\R�@,'y��N���=���p���^Ő;Si!���0�G�*i�|�������x���S�)�H�ǌ}�X�����7�״Z=>��Q<V�!�m�}�p��A!��)8)�ڃ<N�1�҉m]�7"K���vZ��ĉ�)�J��4CR�QMқ�n✙�u�b����ϖ^XJG|z��A�
�MF�F��,�}��s]Ä�S�Ѥ�un�sZ�le�\��}�`shI����qh�C;V��a��������<��<Y��E�F%;��i8϶��[5m ���9�4�n��ٓۉ+�>-�	�V굩�d:R�q睈��X��OR<���'�9ϣ7X3cm�9���z@yv7\!�qutu��󍞩�%pvxu��%س��dmG==�fK����x�μ^�ңQE���\֊�[�shۛk�W���!�y��E���lV������0��
#��P���x������<S;��b"|F 
v��N+���>$�J_wrs�����F)M�;�S�,|8�ڇ��S0kc~���d������o��b���`cD��r"���l͑��ӞxO�$���P���c�-��v�-loej�Bb��˦�N8P�f63U`�qȭ��N����xJ�ey~r#�V���#�[��"�TkZ*���*�;��t��!��
R���r�%�ns�kUh"{�g�Dq�����XR��,3Ԑ�J��W>�����<ؔ�qZ�e-�4fQ�a�e�
'�6an��{
��iR)���62ҮA�������Tp� �bW'g>�E�V���+"1�>ۉ(�F�}���:0�D,������ ͙��M	G0�������W}��ͯJ��sb�ȱ�̅D* TB��"TgV\�wzחw8'J��s��D���񼣌s%Bj�G�e7��N �����&�vZ"GJ�Fī�m7gL�)�T�ߴ|_���u��OW�cDC�8���D�B'��<�Qi�D��4/�u%��m�/�-����Dᅰ��m��m�
���J%�}�l�P�+U2I-EX�v�z
��볣]�w��}�\���j�E�D$$dRD�B���U��efK�Sm-�qւ'v�N�A A.=p����r��=Z�v5b��ˀS0j�+�43�nj	�A��F�>"�<ab��q7��$7���
���Fc�94�G����*��p>�x�>��8n��ߟe=��7x�U�Ot"x�^�5��Q�v=�3k�3(n�y˱d�����ic/�d��&��h�wBTOP!� �qQl[��1Ix��j�1�]�`W#�+j�if����Yӯ�]Z�3Gc�6��zORv��tҋ�$�WU�Z���2퓕p�f,���لա3�ˢY]vu��a�����M�b5�[�������/��{�1�u�l\���00Xih2Z,*g�
h#���	�8�׃��-�2Ot��R:b�.x�QA0��{��>L7��P6ʎ	0�����&L�R>�'2]�jG�q���߾V��<abV>�r�m���l��x[O�е�P�l6JHѼAt�߾jij�f"Q
����v�+�oa��,�]���R�}�J�K�93m����3�����|/�]�ε�T$U�Ci#F
hH.�0玨r�τrN���1J0fo��qE����}��:�����$�;��ev�t�����S�V�8늭��V��g�
Ń�	n�g��ϻ{��n��ϜlYD���83{�}�0\��̿���N��[��S�#QG�U�r۫�?=ʻ��I��_����>��n�c�G ��id͓��*   �lsEE�X�A�޽�x��O�n��g�E��c|mF��g*�)qd�1�}V��4���5�p�&j6�6�#]\9��NTn���l�&�|��������f��������) !��sc-c���Q��a�'�J&���h�"�&}��� �R��o]>Y���]��엋�j�cV�0_T���0�����;���Z���s��`D��F!�>T����*8$�3ڗ|>�(�_gO'9~w�Z�u��&��H��r�.�T�gAK���}��	�|ݍ���))���|L�y��«:A�iD$�WC����st�<"�"'> ���.=q�|g�j�0т�>����L7�=dUl	Ț���q���Qѝ6�.qNuC����y˲����w'筵����s��v��=l �5k+����X���/mNu�JnA�Ԗ�hō�"-�B����>`��SZ�c�p��Ƕ���5�`�^`�j�]j��=�~N��{���/{���}Aad���uVt�R����V@�{mͣ|�~}&�>��)�b��CD��_ug�+4g�iیgO`��@��Vt;���+���
p}�dр	��t�(C15q�yoM�������$�m�%Cx�:�[�.`�j�P2��ߴ�1�Os�7X��ϰ=���t⪚e�i2��N>���Ӏ���̭u3˜�̵ET����+(MY�>//w9��h�6(�+�ݮ��ŔM��O`����a�0����7��8���a�XhNi��y�d�����&g��&w���q^�߇�����_XZ�e�..p��|$��[�֪֒.ر�O���*�43�n�:�*b��|"ՔO�V>{���D�I�A�o�3|�w�Znh�s'bO�����C�T��N��f�C��,���J7\�X�p��S��a�jʏ{ʨ��<r5���e�H�Z�U��	��Y3P3�wTm(k�Ua�o�Ț��7^�[�=i<���fb��s�UV�V�#yFv�.���_�.������)�=���(Ʀ��ޖ�Q��W¿8*�h��&H�����;&L���`!=Uu@��*��Ġ�:^�إ���մ!����n�c`e��]��Wyf������wl2gA�
��y}aZF�LU^��h����GQ4Q�����&lS�v�p;P]ZQY�X�k6�9�(s��r�0K8c��h7��=\Bw3DT[�9�ͽ��H����j���Y�st�W��j�iNn�2%�&z��qY?iW:s\�أ�K��:�΍�o	�y]]�YF�*N/iIٍ������i;�RȲ��Wy���a��U	vk�t {��}���Q��Ȕ��m�~�ׅ����>~�징�Qv�����x��#���/��<�������Ѽ(1P�wu-��4�B�^g<fe��}Y:&A3�tN� �a�����Ѡ�7�V��y��/�Q�N��Br+��x�vv�+n��b�����=ۚ�3OR����+�F�/v�y������6mܡiP�F����e���;0,�Ok {T��Pq�ɾ�F�s��z�No�|�.�߈���@2��D��w��j�I��OrsDX�jв>��y�7�ybz7$Ʀ ]���&4��� �~��PH2H
�'n75Z�f��0�ϟ|j�A/�_�$��_̅�g={&���Sp���u�F�{o���rJ��;��rY���Az�E��T}�偑�W�5����ʩݘ�MU��e)�n�T�Q�H��me˚:��u�)�G[����=�=#Q���xuԭ{$̒�ӸG��Xx�MF�\���}�#�l��������eIW.���<��GPgT\nx�S}h�P
�/�}E�n��~��xK�Z��Z@��5@�|��X@D|1\�r>^N��Ë�l��[�ٸ������1�e��$GW^wS6hљ;�s��og��:�!Q�TR@���;��u��zs	�ɣq�|�܀T��J��5A�r���!�������qe�MT��5����a�9+{���ԝ��G�a`djwՎ���~	`�T�]�n@*<�K�U��@nr�b@*7}Q���Sp
�k�GQ�W�xU{�XVhu���29 �X[�8����+ �j�F��hߒYXf��P;�y�P
������<��GP�F�+�j:�u���e��N�Os�k �jlH��P���A�� J�_2 ����*�]1/�BJ��kU[)̜��%!`��<�|�o*"���6ozF��w��ɚ���Ȃ��p��7k��Fl���R.mep��E�g:�6+N㨮յ�L�*�Щ�[-͔�u̙��e����.��T@�"ŀhR֮`���S7i��k^��ݡ�SB�I�m�7���	e����8Y/^�#�R��9���.���l!(1�9$��ֽ����yxY���s��wvdj�XY��@�y^r�I����.�z�7�i�9 ���"���RC�nǂ@A���ٕ��֒@9�-ȧU�u��P
�{�!pz���g^�%˽;��"��0���}h,����W����0QiD$�O�#���}X�W��AM���Z�0�

hk�&��k���]���;��&Z"&Ov�V�'���	?�Ċ���? ���h�"���f����؊G���MÛ���cޜ��j.��P��6�,�YP\��2�t@��.7��9	D�h�RT�Rz �7��2'���C��fG�K�xwܭ�&VT�4�Q������wt2<����}��G �e� ����[̩*�٠78�.�Q֨y�٨��p� ��ܰ25
��o
�/.��;��dr/�!M�%��Tw�F����Q�'}��I�P�ɛ�vψ4Ƭ�}6��[���kRh��%h�5 �[�k��b�j�>j-7A��29 ��<�r���SN���ÍA)D�n�:���\�#p���ت\y�~��U��@n5n�F��2937��_�����]�^��+��zU75ن)_d�n%��Z��
�q9�TYɈ@� �}�w^�u ���Z,�B��ҫ�u����w�iD<�,�n�X[�
�C��X���!p�(dn.��'eYXf��P:�fcS�E����j>�펣�9���x�'�rG��}�'��9�#rM�GR��U��s�NY����0�4� ��~K#P��dn���u@7~���\��{/�{���m=%
#�z���27 �-�G��X��7�\���K�������j���N$���F�ιc��]_�~�VJ��n7���4[�G��X��e��B�ٮ���G��XS;j6������3�B���9���v�6>���G�`��!Q��G���Q�����˹.]�;�Tz�#S�`�s�X�;��r̍�:����o�w��eԩ��yxEZ\cf�l�sfi�$�����F�^�=^~~��y��dך�7~�<."������wg���tUhu��fO(&@;�E� ��~�F���c� �q���K乣q��� 9���$ �p�luA��nF��+]ɕ�.�;��������5����Aߴdr' ����[�V�y�*��*�ٽם�fc��~��9l��a���1���.۩��UF�>7��}��B6�K]׽t� jΦ%^�W��]����`�����8���.����i��]��G>�u۞���s��K^(�fY����΍Χ�m�;G[2����C�]��E�'D�yR*RiEx�4HgJ�n`���v�ۮ�T7V���:�r���%�	�y�K���и,�з4�B��"�9��3z��M+������Y!籚��h��[5C��n��>�d��IUeV����rx�;�r�I��C o�80 7�u�J��Zw�Z���A򻴨[�܊s}z^�*���X�P��-��).��n@;)���$5�u�U̺��Л��rY�j/�;�E��T}�偑�םX��ڜ���TK�%�F�Vc���N\V��w����Նh�:�r������`djo�y�P�Q�W,����9�R�]��?yi@/fHu�B0\ӗ�*�y����a�_1���j��\n��\"�ιwWS��7��޼[�{'�ё���nC� �q�u��L�xe�q�y�luA�wfF��W��[��/�k��V�S���yy����(�F���_%����k��M��E�w���u��ۻ��K��n7��nE��G��Y��^�����Q�ȽOW�z�g����e�.��+-n��h;(�;y9�Ni���ԭ[�z��^���F�����u����J#��^��܀Tz���s.ꮦ��j�-<H��|�Q�W� o���p��y%��R�u��#d4����E@v�����fO���ص���k�� #xS�Ә��U@�Ϣ�����^�9ܞ����[���AZ�/r�#P�ucq�3��P�ܹ�q�F*��e��Tw�F��9�>�vj7 ��ɫ�L��F��*>�%����E�ucq�C�h�u ��-�G���K际�ۙ.	�4%%!A�29�rNvn�vi��f��5=�����25 ��B�Cp�/R���+��s�ɗ%���w�h��U��h� �����w��yw��vM�̒��Z7�s�[�
�WԵ�E�n�F����h��W�+/*����� ���F��P�r�]���^�����,�t��p��|����'9��Һ�����4^���a�ؔwխ__o{��U����ˣf^�@n5
�p=^�B�]��@7~�rQ��25����_OҌ,�7KaIv���+b��z��9��w&/g7���]�l}^�� W����W�\v��q.QS7�����̯:��L҂9:7�"BHM�/l0���Z��G @u�h�r��[�
��<�y*��h���:�A�fF����� �y��F���+�=.��ՍGp{���E�����@*;����;�.G �O;��u���z�W�-��ï	�R(�t��1;�#2���Ү����M����4��������VzB���H%6������q��a��}�#�T�ܞ^���v�����Wf�5�v�yx����n]]2�^�فB�3n݉�Ri	T��<M�ٜ��m�T¦/2$Od��em�s�%P�M�����!�i"�,��VFƭ��E����r|iȏ�=���Q���@q�*R���)�8[�ܧBM	��\Cuc�8�~::��=u�.4�E����`�"�{�|��t�=��K����\	�<ݵh�e^7�iS#FF��'�eOQ<�Owu���|YV<�}z����,'[�H����$��]O���akRZF�|�{������۞&�Β��pb����@��DZ���v+Y�ϞjD�WV$�㼜��JuF.	<�UD��
Kf^��
��V�Ж`�Y�����
]c�BJ��c�o4�4��F.1.��,meV�"F��Kx��54�vΩ��Ǖ#!���*��7����3��웵��v��^��2�c����k�]\�4��aI�wl�p�BƎ<�ϳf�F?p��[�꧉Tn��3>\�������jw�"����;�؎��{<�.!��j�������cƽ�u�1(��Efm�!�q`��w!��F2p�@CZ�]��0r��p�+�`�6���f6K10x��a�ֳ48H򕕚;gC9�ر\�+D�Ĵs�X.֘�(�n�iu��F�%��r�����a\�y�
霮c�{��H�uF[8�hV9䃨U��Y�c�1P�a��>�<l�mq����㗰v�n�ݮս�%��5n(��eꍋ]�>|��?2��lp<ێ:�ĩGg[��;(jݼ�.����<�\�d7h���غ��nI\{r���.�r�YV.�z���y�u�.��j�vŮd���s�Q<��nJ.�����mw/��B����7�����N���-z��A_��(�"�ȓ���n�u��;�6ˢ�SɓՌ�e�v-�m���V �����ьC����پH,��WN�Fk@5�&���9N�<,�'n�O~����Sv��$Wh�[�Gd'�Ӝ�Փpcr=x�	�{���s {��q���T��d�s����x.��r���{���F��b��8(�tx ��ǫ�7�s�=�԰w3��ݴ�ضZ�����B��z�fᄩ��ݗ�k+�L��p��>^�=�=�o���5�p?P��g���K�^p�'�P�(dk�/
��zk�_���wW�\X=�CC>��	�dd�ag��c�\�v��J"�7>:��m��X"6Aq�'Z=~�^C6RCe��iH��Zۈ.*�A�][�##�l�����e[���5�{8K��ȇ����׵�@�0������v���<�D[�,���b˂Q
����;99$��G��!��j�[�
�W�U�j5��~ AQ.j^Q��G_f˩r�ӹQdz�!Q�w��A�˳#Por㾎��J�wUwu�7�/��A�tdrpH��E��Tw�F�ݞ�%�u��G|;���<՛�@:�r!D}�uX��"�\;�lj9y���K�7�:�rS����U�_	�y��������m���TyNM�\��g[�g[���Z��T�*�:������깕��h�(�:�o�-�Gg<�W�r��?A�|/<DǮo���İ��J��t�	Z?n�i��Fػ	�&1�u��U����"T�T	=U.5yvdj�0� ���� ��+��'��WR�YycQ�{FG �r' �!�N#v�>B<181Ċ A@�{�u ��|�`�C��ƣ�����Q�}O+^�0��i���y`djp#�(uA꨸�5�� ��''����鳶�I���bu��sLM����ν�`M3�c�OT�~�eo���C^�g�5 �אּ25
�J�e֍^�u��=�H� 뽖������5�W���u��L*�V�q���[�
�����|=X���v_6��ȟ8Ķ�Q��nO7�a�wg4@Q ��	$��q�k�\�A�Qp*���uWuXU��FǙ﵀j5���Aߴdr%' �ߴ�)�G�̪��2����Зċ����{�rQ���a'o>s����[�8�Zj.sy�1�@�5��M���rof]�8^z��h��Wܷ o,��]F��(|���qq��2¨������	s�1�� �zĞ��F"��?f��Fc3���:�#qw��"�|�޽�2���@nqb�9��Tr'\�#�k^լ��y�}��B�QJ����Z���-W�q:zo^r�{'MюMˊ�\�y�B�D�j7����;��d��wwE����7��Q����F���cQ�<��%Q���V�/ɰ�s��g	q4�|&Hq0I@Ȳ,� ,�G�@~��L�C�h8�]GPgT\n��9}�j�;�T|�=�D��T���ycQ���#�
׵nC� ��aUæ�]�w����r��F.���@�#y�{�i'o�σ�e+���y���
s�5@+|�rQ����t�n�Q�;�'����U�h�n�x[�
�'y�V��;�lj9~Q��W$P��˻�2�v�Qk��'�DA�M@W�����S��oWVp������UԍJ9v-�.s)�T�nh�ۛ�Ci;n����`&����2��a�f]�E�[�?��^�
T�칗F3��i��"$�jp0�#M��ӵ�m�+����dGk��o�-�%�aS������P�A��-8�1����ڧ{�����<�B����dj�C�ȳt|�ox[�
�������*����5_��`7A�kT�^�V�S}]�H�5�w�%W2�U����]^��gi �s�kA��#9�tU�a':u�z%��n#���q7���#Q7��{+*^�=�:�OA�}�cq���̭{Y�Qz�~RvْhA&���k�,(nl���J���Gj�I����sG ꨸�ZË��q��,�Cβ#����D}�@f#Ltol�,.��l�F��F(#��b�Nz�}�h��9���:�:��0@��~�E��dZ�n@+��dj�X1�|W��Z2(�;� �j�~ ����ln!�~lߦ�]ʕZC�`�̀�H�� � �az�g�����;�ۏ�{�Z�^��d��!}Or�ֺZ�:�"	���s��MٻS�������߼����|&�
�=�Ԍ�����������Ռ�!Og��P���F�)�8��W]��F�6{jރ�Gh�#z�s�9έꉒ��y;�9�!!E	�
qs���",g�(�� �p�+�G�d��ԣ̥	��{�����YU�ܓ�zV�͡�It��f�,I��]�.�ȏ�9���M������:O|���>����ؿ2�a3^��Nb�Y`  ��Ĝ$�)����}���
�F"ډjV ���y~Ss"�O(��=�9:�2�pDɽyp�]�~���椂n# !�מٓ��A'M{W�����{�OE��n�8!��8�b�T�\X�e�A�i���0�A�bS��eW��>�:��3
o���#�7�L:���;qQBrA���C �Jo5�#�ͥ5]���sk�K���]B�1��0*��8�#ﯹ1�Y�;����lmJ,z^i��̾�-�gU�?G�/��R��-��z�72�.��9K��.�4����Ě��;wN�l��s�@q[�����u��<A˸��&69F(h�U����^�sz���!��4y���״�y�#`��˝��hʹ2��I�/%�Kd嗒f�Ru�5MiK��hL�GYM�����f���=�������Z��5SԜ�(A���}д|o��(Ƥj��8��k�7�X��)� ~�ޙ΄L�-�� �4dg�HH�U|���?Q�w7�}�/���O�Me��ғ6�,2�j8�å���&��`���;�������@�čz�g�&h*�
tPg�}�.ⳑqj��ۖ��q���䛩͵ll�}��b*qw O����Ā<>�[13|��W�yC�A�z��l6b�7����L���>�M��Xn'�i'�Z ��},��mϛx> �\����kP��F$���>V�5�쉘�� ��Ii)��CD����4�m��)0����{�E8a�u����a�����#�*�UB���a0[Q�މ�����1Ë�n|���X�aBa�U�L�ZP=Yy�a�#^��(\{{K�g)�O�[ �X�~ۨ���b[���$�]�z��ez��pw3F�/T�����e�Y�ū�=�����n��uP8���8l�1�c1�ofm�Z��27�Vr���u��L����_Jd�\�㼫����43���R�u�WFST�8Q�&�݆:?Q��먑��y�v���%B�,��y,����m��J���o�����͸9ۚ ��~�l�M�s�W~�mm-�ʮs]�ڸ�.?m6je���=���C��m��xw�{~pb��Q`���k5dR�y{�Y}���MR��iS�p�9���[x5�������4�|���8?S���]f������4����:?>�[-��Ήj;0geZ�llu��͗�J�;0��2����D@屮4�fe�7'l�?:�?T�K3Fq����p�M/�M��v=�?q�>^�|'�q�vرi�xk������}2�k��U����Z�P+:��R�{1cƽ1
ɹ�Y2Gm����Ð/��9�'��qZ�~3�篼=���٢��g�zߐ���1�G'��w�W��8=�3
���6��n�M�,���N�<�wh���{��4�P��G��o�55#.���/,Sv�I���*=���� X��?P���9NK�Q ���V��/^������Ɗv�L6)�Ze����s�
̂ƶ�@.�H�/\���^�Ǹ����a�u��,ֳP�0n,[��Eyl����Y��|���Fq���'#��Ə���\O4�~����!��M�+��ϧlݗZ��>���x�n1in.����n�� }�L���M0�f>�}���sx�4�J��Xn;�1q�;�{���V�e�B�6��
J���7.*�fo R�D��������@n&�n:Ǻ��A���>��S���n&�v8���{Ñ�EMG$�0� @Z�[��p���1#SZ>?�ˉ��3�L�FMgޞ���;��� �+�_OY�ŁŪ4c&u]�Kt�WG| ����ER4.<ʆ
�ž����}��L_�q>��=���}��矻��$�jQ��u�!0Q����	�\�Z)	��l���)���0$�[�3�5(G��SQQ�~q�H]�7�7]:�UE��a2ȁF��n-fD���>�?J��m��+��ˈ�ߏ�,�����f&[ �܉q]�����QU<ӎ����ˊ�7L7T������M��Y�ӫϴ�;��<c����	��{�_~�kO4�WX�f�����˅+�8E�4��ڵ��_�������̐��ۣk��;Qu�н� ��]qå�RѬˁ�=T�8���x��9�aM�ZW��r^�]�".�3(��ʻ��,�Ȅ�r<O6ʄi���\U�ƌ��e��L?�;;���N������w�~	?W��4��l�:u�|��܆�=~S0i`�?�5B���a0�����D�ָI�Kq^�r��m�
e
�}��j���+^�L�aCQT̪9�[-ݰ�F֩�������lk6���\U�X�%(�hv�9(˜�1�z��M�ș�~|>�>�y;�>�%*�1�o{=:-�j2_��$���;��gOov<R~�6�x�xw���hh�C��3BD�)PI<�{��Ur�xgHj���l8PT�;����	�����G�#�T$��D�M��yx�}D5}I��=��ME���]Ъ�g�f*}�vz�[�t����n�fmv�F��W����ֺ;\h�߳����yq���>���CqCx�:IiBQ���歹�*m��W� e�ġ"-R���q9��z�C�˫��x�cR5��ȞP�ɈNaT;qz�V]5s]�@��ϪzT��]��#� 	�~��a���)��B0�a2�Q���BfV<2�ߚw�s�v����."�V�q?����Eo4���G����Gl�K[�l.�6�\��.�`hg�w{:�WJ��/�4����p*����"5�mT�\-��q7"f9x��7�~��;�u��u5�n.�{�W��3��[_������8�zf}]Vҿ��]=� �i҈�,F��[�ݟ
މ�
�ӡr�� '�I�˅���P�(UGg�f<>Љ�oc�8,�^���X� �Sq�חXxe79ִ֪=c�jĹVw޹���⩎�"��m�E�󆁃F��>	+^p}�8��߾����i�Pb*�u���J�em��G�{���@����31~���"\�F��T�\"�}�"f9x�����x��ds��qb��:3�k�3-����+c�r�K.S_s���Dph���k��[�����Y6p=5�i������J����A�0�w<��8S%h�<MO�^��l0M��^j뗚m�Z�� �mq��
v�j�1:,����-M����9O���8��s"�0ōŚ"aTi�;��o�7L7O��2�c5�#e��9x��Eʍ�q�����=��LW�hh-(B�=���G~�"\j��ش�"��b+~{�U1��Sx>m��1����^����+TTyÎ��������+2�Y75nkG9�,!��s��vLk�A����> ᭹1^�
M�L��2<�zU���Qcc����(tR�"x�-����wLdUvmd�QyԱ�	�]"(�5��>��,�H!	��Z�w�fW[�8:��{��j���E]0����詌�8pz�@�Xn��|z&c-����y��ReO��|XL*��z&b�Φ�f�fb��'����v����-R3ൌ�n`YA��-��Q�g�g�c����>ڦ��L�b�<M�Tf�|���硸�a��< L����^��Y�7�g���y�u͋��D�W�q�uN+�j&���ç���+۾�S#zEY��d}� >�
��qy�3��i#U� ��K���T"��"f=~3�8pRQUp��^mUE�������_W�֡͠Xb��0��3r��m.�Q��G���4���� 
��8��#
��5�}�Y!��6�_��;&�A��A@��]虋�q�	W����Cq<n��Z)
����qp��0���M�{NXs�rM?Tl�L:�����LN�s|��\X�� 	�|	Q62��r:#�Bu)������.ș�����g�@s�8�"�'��!u6hQ�Lm�L�,0�Qs��qk2&b�Ͼ�b����CM2\I�C~�e�FJ
���p�؄�J$�qSV� #��Aձn!�8 �F�v7�<��Coe��O\#�M�Ͻ�у�*��Y����T�3�˧�	FO�q��D֛�ws;��^��9���+�w�:�����1_=Dt���j垊]������>�fE������mE�%==;�V��o��>+�����%�Зڽ�˕3a����LGA���N(UDO���ǚ��R���;-�?a��x�n���6:������V!����E�)�мQa�+͓�{KY�IV����4�o��xoI��f�<��5��c�w�!	k'�������_Q� �<|�ٴ[�si�S�'����}劷po���I�w�q��<6P}˖pf����q:�]��2�c$���5Cq(�-k�,{��G��ǣ��r7y^�UX�Ӻ��:#����5d���Q�`^d��y��j��E(r;'*Fqp�͢����cv��|����t,Am�qAA��r�S�|֑�.�~��Ϝ��H<Ks�e�dz�����r�C��v��Xo\Vޛ�n'��Oz�@��ݍ� ��<S�iR<�s�3���-��MTd7���sc��q�1 ;�����c�,i`�3@Fh�jF��1�v���n��c��pS�5�b��q�%Q�1���Vl�cp���gc�M6SWeɚ,����P�2]��s>�gkgrV����A�2�7HM��	S
XCX�kc(1��.)4#��xٲE�eZ	�x�7m&�rݴ	1JA�j�48BDc+��%��M���`�l�H��da-��ѱ���),�B�)���6�t�ָ��j��+�}�,G��Q��h��ډ����pq���Av�l�u��]�����ps���K��/0n�	2+�^�#H���s�PEm8�=�1�箸�<�)q�O7���hzbͧ��Z�z%��#g��;p��s�4v�����c���K1	��4u���9��kʷ6�.u�gj�Q�ݢ�8���y��4N���;��W��+w�b&5\Sp`�م֊gϫ��D��P�#J�|�Y�%p��Y����������G�H~��w�!Mw����c�=G�.Qɜ��q�Hً�Uq�XKJF7���&p{�K~d�@l8���9^'��|�����pdrs�� �D+����'a�}��=�g�&n�7������Ջ����zq����9�8�^'@�������7�o5<��d�qi�M����'ø�vY�Y�,]�S�y�6�0�KL!��aC�<��~�r�GцL��뮇��4|a�G�5Ei�-o�d��<���F��y�B�n��^'HGu8D3p %M{q��b�����#��Z|�]���3�W��㓏�h %�#���	d�;"��Ot��3��.��n�j����f��r��X����b�k��m��O"Y�1��H;����9���6�k:���+j�aFE�l�{p<]u�)rq�Y��U��2��+.��@�D�I��yeo�V�ҙ�b�� a0Ri�`��,6AbN��2k!Mo��O:����/E]^f���dI�G��6`����Ճ�~����zfb���څ�h#֔�FR�p̜�5��5а|*�gs	E��"Mb��3&l��A�z'P0Y(���i�m]m�zp�]��r��s�)�l�F����#����sXb�3���eZ��.����)¸��HE␎��?�Q��(��~���nw�z}�Hq�v\��\�߈^rJ�]WwU'�t�}�:ң�i�(v@	oB&�V7��gI���-��Ľ�i��a���n0A�k�/}p��1����p���wi�E����ǻ�3p�M����
��ۋ�8��(5F��>�K2�~i��߄��T�d�������Y�K#]*ۗ6)�R��fͰ�!�Rpt-O��_�֯\��y�D��! �HȂ@$}���+���}z)&a2b*�|�zS�͙���{��VH����!����V���hL�w�7��>�>&'BPJ@�&�ym���\���\V3�����q6�q�|>�W�������TGz|8���G�m�Tg��P�\ ��*�w�7K��ʹgy��B x4ە���}1����qG��k���U��vr���7�	��rof)E͹� rQ�|�[��]M��$�I�E�3�Lz7�	{�ѫ����y���+����'=���?L��A��K69�9�mGe�雕ף��6=z�������{�a���A�>�+3ff=��M���Q�:2��+��!M����ř�n��q�F5DC� o�f�}^o~E���A��AEVr�D���Ι7�n�m��"s&����b}��UR�O��=6(Г��q}�(�E��y
����. ��"�FGBE�)��4�%�Վ1ɠ�vH"�݀{zN5c7\kc�-�F��5.��:9�����q���6at'j[��N�Jܴ;��Kb��΅+� ��v�=i.��'���ww����� $�Dj)y�U�UcYum���ț���E�ց�֐.E6<w5�p!N��'����1����j����	��n�Q�ӿ|4ݼ�1�x(-DQ��Ŭț~����3=c�0R�J�����9��� d�o���&mI�� ^��{�A��'�'�S��F�ś���3�S��Rm�pd����!��o������cfc�De��U�\��BP%o��$��k"3�cN��I�.wn�V��y���]vV���)"�!Ｒ��f/�}zϻ��`��G����	��7^���&!N��B�=>�@[ӝ�� x4��{�ﾝ�7���~�|MZ���kKǓ������P�!'�o��S��ָ|gK���J"$����	�h�%������.,�EER�&\]㓗�9w :
� >�p��	OY��f�v	�O	ި��{n!\���ͻ�w;+z��{�~��H�� }�'�>Ѯ���@ر�B��,L��k�ż��y�Eǣ댃�!�{!��r&c�ј�:��ZA��G����kr=�\�۝{8AE�G�5���g��Lױ��r�I�.@��G���qX�U��"�M�t}�nv�=��l3ݏf.8��與
��i�U��p��ԣ���~d��Uױ����JB̂���' �Ny�sz���\!d@}�^kZ띓�KV�L�ݹ�}�ͳ

z�l��;.?_���$�[TgƺI���(HB"E�\&���g/�_ &r�F����7��]c}(��|&�b��nw���~G��0!zr7�a�]V 9x�7��_��{&n�r�'	�����~��[�3݊i������<y��r��v����,�qj�Oh��]�&`==�����;q���J�\���m�vQu���n{fB�l[Kdr�=���S9y#<T ����l!�eN����L����[�)l�q7Fɫ�h٫h��"�e/(�˜�RFAR@C������F�<����O���!f�;)�&�$ڳg��������F�P����l^����^�|�{�fy�};��]�|"�IDETb	ESy��UC+-���+ŘiBJ����PN+6fc���*a���c(U5���1�S0}�8߾-�#>��b(�Yͻv�\Mk��������t7�Q�c�~���"�_��J ����;�ނ�B�c�j1(c�n��Ո9,!L�g�ط��e��̜��WJ*���+����������x����`I��q0���~��3����b�zl¥Z ^�ULv�q(%�.���L�>�Q�k� �"f��}=��{��ߺ����h�mv��]M��+����.qQrP����<���|YV�P��(B%�J��9����nl�ǲ�A`��ϲb#Cj�!����8`���V��������.��2���?��F=���y&<�r�����	��r����z���9{�$�Ѷ�ުq�T�l�w����}m�!�'��
�ѱ�y�b��59{u�Wv�P�c���*~�������o�|�]���m�;2�)/F�"�k����f��Þ��8���G���v����d�*��,�L�أ����}�ol�V�е�r���wf���/dm!�ԉ�<	��ƶ���oo����޻q��<��DQ�̍s�c�6޻\s���^�O�Nn���6a�=��{/���s`�8O1�;{�_6��%�Y�4���1N��.)Е]��V3bb{+8���N�a/���6 U�� �bo��^6>>L�9j�5��?�<�������/�|�T���x�jd۟	���e|���A=�!\�� ��f'�1�@l�����^s&�0x��@����gy6w�}
�a�ߙf!E�W�x���{�w)�E���Q�,$׸��>�o�=O�+�ke��q��g�DI�Ǫv�o'D
����s�H��V�:�ܑ��p�QSq{�^��y<��u9�x������e1�<��)<�O���0s�F�#���88�p�2�f>�Fiu�,�Ab1��<"�%��4w��Dч;S��-bJL�����Z�Ѕ+�u�Y��u6��
6E[�ʙ7��ܯR<�L�v�ii�v��t|B�����8�gtC~{��8vnC��9��^4�7NZ���C�v�eZ��8��ڈ>�
>��Nn!���7�<;��ldW;*YU�+��� "�}W�S�e�K܈����ﯶ&b�J=M��*L��a����TF�� E쩏g�f=p�o�
����S����Y�0�KJ�70��t*��^��v�F���y'd�B7{y�ڪ>�x�s����X�*���^��"}��U�߇ҍ�S�Ι��>A��"��ݬCk1�P!z�)�tV�Q�'/疛��@�[��@�"on{n�R��.`6�z�]���g��?���~�\��;�q%F�͝��������t��9�օ
{/؍K4t,.8ўx-R��n	�qv��ι��E]0�F�;��U����B^Qsq�sG֑����>�(p�����7���>�=S1Wpp�BwﾏsF�G������i1�|Hl�Ts�p�^ڙ�c�cn&�=�/{�;1Bi�P��6���S�R�nul���v7�);cYk�R���X2�q�6XY.�@����A�5�*�����;�tY�Z�\<7=sD�զ��=7t��R���;v�=&Зl����p���;S���ah*�y3/(��e�^!���! 2,��wppy�l!����)�N)ۏ,\��%��lqzI���[�./���Wͽ����K������%fKqp��a�Uo��L�CP*�|ۊ̙߀��Jb/n{�F8���#�����\, E�D׺6�}���:�})�X�w� !���j̑x�o��eƦ�2�p��Gl7���{�ꪏd7c9P���T{_�7���4���u[�&-Y�P��1�ydI�j3e���7쵎������*H
HH���՗��[��U{�Q�R�����f6���L5m��Z+�1�o�kl��>�X�]��<#���*� ]6\������A�y+Fz�B�
��n���of���`��-�	Ey#5m�8	�T�Q讄�(P�j.a )�	F��L�y��e\�-QSQ���P[wK�J�~�GF[1Ȩ�#e\�f�b`-��ɶ7^k����Y��D���$$	:��֕�+�p���(Y�����E�Fkπ���YȆ��с'֑������Ҝz�'�χ��$���(Ը���F��t�1��쾷�����O6�C����li��TQ�K~�ڲ����g���BP�����W�	��@j�xL�8&|}軵��_�xifnġ���2nQІ�n#��e���4�T��ܚ���Z �|>$~ ���|�^�s�n}��
��yU���l{�����\���q���v"M4Jf�Z���r�4w��>����~f����!�˅'�g~+#݋��w���^�a�W8�L��m���f+|5�&��[�K����Y�� =m��"��M�`���⏹#=m�q��P�,��鴘*�}׎+o�F;����g�"D�xFRU��Q��(���~��޲����Whu���m�Z��*������[�pO\v�mNz�Ս����4�gq��9���{v(3�ͻ0\��]�yNM�9[�k�`�ݦ�c�7��Z1�u~;�������x<���|��-A���{nF-L�,ū�9�l���@�����E�x ]D?Pcd�Q'�[�32f}�n���}	-P�]��B�］Q'�#0&5��a�����f�q�i���t���#5D8J�����#��fO�[��{��}��6"	 �.(b����t��D+k�7K�g���]�� J�Qf�LG���Ts��5`�k<ǳ�"懱���WGN�o:�Cs��4�ފ��ٱ�י�C+�F�1�-*�67�o7t�>��>qQ��(<F�D�*��7��oj��8I��W|k��f|�π���"C���'�k���W�>��n����=y�����MFa5�S&�^�T�n �OR�������#��#�[��4�mßv� M[��ٟ,���[.*�Q�N�<3�(���7(�jkʨO9[/�e#�X��Q;i���U
�<�j��A|~$� O��I@$�O��n{[���D�'�G{����}�\�x(�(��^�wחu��Q�H�)! ��am�,	JM��m�b��ᨭ7N_t
��Y�v�"�QW��ᛌ:�;���ƾ��Q=ц�D|��U|�7�	dC�S�|s<��57Y�O�'nLq9ha��������\ƒo��	�Ңcj]��7����	���'�H�0�$�d$c	���+�ug�%k;W�Z��Bg��:OF�,.ĳ;��̰���;�v���p�^�sۀ����Ŷr#��ZP����>5Z����
���>p�gy^Z�W�_!3����EDN�7�.����յ`��I��;���z�וLB�PF��m�v
ˬ���XD��
��/e��l�10�^W�6�]�XY��N�<A��-y��ں��z�[�}��ÃPG _9P��g�F�S'x����&�٩R���(q��B����{#.�ȿ�K��;U��d�s�����}�b���-�>��<�9B�}H��Ж�$�r��$}��~]��`P>����fס{m���Wg���)�JЬ��ܴ�&�d�4��<�~�?�߬j�"t��\h�r<��z����;����^3��֑#`�u^��Ź&^U�v&����k�SSP ��4�o���Em��ɶ���p%�Vh޻ݔY��48q^��L�UڟTN@�Zw3h���}�wGv(&��[n���7�UoL)���{��d��ﮰ�ȎBX	
��6Or�@�Oz��-�GJ7CO'V贳��+�i�r�����g�_�W�Ca��e���!lʱ��X�J���Y���-x��m����ڇ+�Ja���32�u΢�I�r�Nm��j���+n����$�u9�gv��q���R���lg.�bu亜EH�-Da4������籴���"�b{:wYj��^{�r�왅K%^
捵�����3��4l�\��+l�jm�CV l�޸��´L]��K5�M��5�s�LJsn��؎�X}W��W#�M���Χ���v�v;zL.����ޣƆ3��Xo-�➩�k5�筜�&C�=Aiuݵ���nVy�����q�b���\�j�j�U]31
�)3GY]/4�cn�n�ͺ|���yϞ�b��ڝ�\�Gu�<�Խ��p[o5���[����b����cW�|z��rEmJ�l#����5h5e�7­�:��IM	.�
ۮ%UY��m4^����YX�JjĘ�@��MKm�t�ݛ��t����3�k�kh��6�鹴����霵40��bP��N��;�͝�BqK�:豧(㺋v�{r,�%LμcP"��C���^��8I@��<���c[7/�,�e`��s�m#9�Xc�x��n�'#^���bM75'N��@8ωP~�Tk�zՑ��E7&��Ň(�K�8}�'*�;Q��4�0��c �#ӕ>��־�����r�4�T�Y�1��/�0 M�M'�n��v�c7��D�ub�b������Yx>�,.�mܓpa^â6�'�q�9�fRi�d�8�3����~w!	��Ƞx��Y&������d�cB$$a$���K�pee�4�Qnc��������~�I_n�b�99@V�N���Ź��ǵM^zlU��gu,��	ø���p![��4^�~Q�'A����O�q��L\tMm
�Ec"V�q�@��M��XA�C	��/3a!3����Bp�d M�@��ղ�̩,�pt��#L�ٹrGM����XV���5R.cg�-�v�M�cKkv۠O-��z�tѪ��4٦my'e��-�^s賳���U���v1q�Ebۮ����4a�l�i�U�ݬ���r���6�e���'Զb��ׅ���}�{7l*�����q�h�3F�~=���G����雼�Ai�BI��}��ueX��_�l�d�K%6����ۆ6�SZ֪ݚ(��YY�t�|>q�͚��"��Q��|8+�>���nf阃og.���Q�N&LMH�rw��Q��]�#k�'S�6��tDRP�J���y���>�`&j��|�I��A�z>k�ݤ���ʈ���&�z����D���	lC�UEb�}�M�T#�����^�&R�i����a]ˢ�i!$��^�7t�>�?}��Ǌ�V#8�h�d.��h����= Oi؉GAh�$��٨Ø���s":��dEo.�T�u_E�s��
��u��9�f�m*މ��^����ǟoM ��������Fz��/��U]��=ޗ���%������ϐ�E���%�P�Z�m�|��~���i�:�Yd�I�����\�iW*ܪ�����][��}�>��VxP�pD�ţ����y����"�o�kQr�Q��SIh=P��/
�e�N'>��T�w[x�(~w�Y,��fH�XS��:�Z*p�y�o,�LUof��R��:�v�+�����Ji�ۼ�}�}>�{w{
��!���_��K URCa�V�q���T:^P�ֶ`$���G��5Tր;P�N_��2�Q��}��J�#��8��R+�8e�J�JϾ������fh�U� ��Z�)��ۚ��*�Ď����s���G�X|�޵���xJ�z���l�i==X�B���bD��doC<�{翳旵-m� �j���[���nð[�|��G�C���[]��G]i3qڅ��d7[+\lnu��	#�ҜI���Om�ۚ�6��([\=��=�k=�q<�v�����S�;gt���8��M��D�w��T��2R��i����2�v�:�pb?�������;~�L|��裪C sط��G�#1����+��
�ѥ��~�W?7���2 ��CE)��{Z5W�+�᪋�Ti��AnQ��~�έ9i��|QzG�qʹ�^s$M�a3�m�=�h�"XE��W�+�(�-� ko[���	CIB��Kޡ�ـ���gң�#;�����n8���A�̗£l=V��]�^s���ʼw@��D��(�|����ޞ>|��_��_x)��0d��5V��'ݲ��5C|c �U������IW������\$�Ͻ���RGԑ����d{z"!�!5Z���	@%W.�7 ��=Q�H����Ͻ����"N�b�+֖ĕ`q�W�*��p�w����χ_{[�ń��蹼���%�83n%ݭ��C{�0J�$W.��e���{��lED��� �����Eg�Fx�mڢϭ*��{.�}�`8$�U�}����]I_'9��~2��ݦ���ȌuE�҈8E�\!75�{[5x�_��&j �k�K8UG���|�G��;*��=t�Q��g���߇��h�qZ'�/��V����v�8��m;���`�Qˮ.���L!� �T��M'jueY:Y��Y+j�� O�A �	I$@$�B����Y��BO�#��K���% z�o�H�!�a@���<ZۜP��;mmBŲ��=�oo[�C�*1!��X'���>��3}i�Ͼ7d���0��kݭ�|��u�dNx[L�9��h��}~oG�o�f����A*�����>�Gi"i�Wj�-U���O��h&��V3d=�P���5w��,v�*����c�K��ф7�0O`K�d�2e�Mo.��V9^�k�$Ʊ��\*�+(8��lp��Q�.�����ƎӷX�����/m���\UqȦݥ�41Qp8�͝U�I��~�x���ǭ�����z�[X�*K-�ڋ)-��֗sj���{�{���*��V��na���� #q����|�}����PCLB}�I���Cf�:��B19������S ��֥
�p�3q�S�.q_�	�z1�,�
;�G;"i��V�����LV�}ujOhC�B
�
"]��}"�t��Xw03cgػ+6	��y�g`�����w���H$�$�		�Vҩ��|rv�K���N#$P6チjU ÿ����Y�v��0�u��~�{|��g��Ķ�~{ZX��U�OJ���ƵUɰ\]0�d�������F{蝜��9�N�h��꺏�k>�1��X�ѩ!x��~S�R�C)��"TyEj�aUK�z*\�v��9Mӳu:)����\ N����W�-���&�J�pmO��=p�1Y.Y�V��-����Dw�W����jܬ�ú��Rq:�0e6$��Њ�tY�Ζ���1%�3ɰ#�i��@�_��N����;oy&-�(�
HY�.�an�ʋ�����\]����S]�.X�~���C���y�� S�o���޹=p��a���v�-{I%ғ�m}�󷹎��}}�WuM}�v#������	=�xB��}v���ͽ���5Gy+=�ߴ�=������H���,-N[6�;�6�ۋq.Yeɫ��;Z�� �ɪ��K߬�p�Y�;�&1�b�=�pX�X��y���q`�{NAqT�պ��ee��V�A9qK�X���9��$����D;��q��u�Ja_�����E�K������6 ��T'z��Ѝ!hj 1i:gdc΅��[����(��GO��ς���í��ۨ�`�nq'���?j��O���*����xr?h�3���`�}Ozzv$9�f���<27�y*Y���˕�"�wf��/�~�,,�	�-��'���n7�̑s���8Ӿ\����0q������]tb�n.a�	-��k8��Ǐ��W��P����9q4���{`�3�nY�kg���j�l�757��u ƹ�����#���(�y��~��Lߍ�oE%m�6`^���o���xs�gc�������NC@��b�&]3,BQY�*" ��sL��pp�G�x�)�V2�6BOڄ�i�}��H H�8��2M��T8P!O����Rx��	�2o�j!\�ϾV�yT��>�b��g�(ݕ�F��d,LOD���]�3)�����wI�9���}����No-�]/��I� FЫ�Ñ���k�_)�����v'Q�j39I�=V^�UC�7|�񷓌�Cȡ����}P6����otpv�:�Kߤb�RF^��y|�wU�;��w�}�K>x�i\&K`G�5���ɱ]��5]�����}v����SY��"ш�ˁ�yj�1C�<���D2�W�@��ˏ���J���3P9�}���H�w�����Z�ƪ�ZN�ǫ�9���y��r��D:������]�s��Ð%�+�$�'�b���t�o�N\��n��+PW���]��21Č�F�=��w�s�7\Y��lkk+��W.,D��ӑ��km�c�<�м�<�Ok,���l�q� ܳ:��CM�raϐ����$��ғ���6�ͦ��A�R-�p9[��SC���k�}�'6o-̈*

Cv��3R�a��Ȉ�AmN�,���J�*�"A�H��Gۯ*2�<�v7�)�1;��_	?O�����=C�x_�2]v�9��C�Sn�a�������W��Wo��u U�c!�l�8���ʲ��mB�kh_A��!0��˴��4L��vYCU��Ķ��U�q�3���?x��ȩ!$�/�\�5M�z�!w����L���t�	��@.� v!'_*f󪱩4`�>�ﾥ��#ZF�������)�4!`�4��fm�`CD6�Bӂ��=�os[�C���RFij0��H�D�4 ��3jn����y��FR���Op47�+�S�J߽���A_X���(�I��z�.��5E��^V�:��"j H� ��H����"�{�Y��4���	�ڕ˩���Y�L��-�n���*�G����L��>�9?N�xO��MG`�̊��9�8z�kCBlO���~����J���*8���s�C^Ļ�"��7��{�۱c`��HI�AqF���/m"��#ѐAn�� /y����]�۞�UK��Y�*�`��D֤�Ԋ��Xv��.��s:K����T�Lu�B6k^"� 	J����]������{��7/U���ނL0�8-�-Uװ�n�3��V�,)*����@=Y'<�i�DD��~���o}�� ���]�1�ዣ��m��[f�>��S)8s`�L堏�0}������U^ĺ�>��_��y���#�9鸞���s���s�F�+#��b�#S˵�j���dö�����4���RX�u��(�5�ڹ�t���2�X�������¦��y[�\���Kz^�qkmq�EiWm�NM��<�8쉫ź+�m�&�g���]A׏Yc[�e7^�[���!Ns�{��'��F�<�<qhM%Y�4���&H� &�&�)����.(������F�_/AH��x}��o1z0 ���	/|ك>�7�����(��u���(81U��'��*���j����.ND뫙�y��Ͼ�� �H�cu���69U������Wd������m�R�>qq�iE#p)����� b�>̿O��L��Q&L�\��W�L�\�=Z�E7�X7e���Y�<��r��n��,�������<�Fs�h�u�h�o�^o;��a��"2���1ezR���a�z�#�J0ڪ=�o�x�$���PG�>'j#�y�\��[vτ�{Z��*UCD1��y����czo9�����z#���R�w��߄b�1�U�uF�&�P""ND�{R�b{U�N{�u�&���S^�i��r��gc�ғ�z��`� 0��?z.[�A�~2DUp&5qYIL+ E('�s�e'{�o�@��go���rz��}�E��)fL4���Цe����˘3#���}��D�{�s���h�-@M$���T�G&��|/��Rquc���{�3}���V0�rFer��6`� /qu�G!�w,��>�*�T��E0��ɑ�]9�q��{v���z�&$��`=I	$d		+[�3|��K2�DU^��}��l�x���}�����A��%cJ�4mm��<�e�f"!	�p`Ѹ�Bi�{���5�#u��y��~��7�u���'"c���}��w��Ao�G�ј�X6����h�G��������.s��ء��	>�G>�VT�Ʉx�v�jVb��]�.^���y�257��v�&�jۊ{��b$�X���.K��y��L>��5_�'�>�(|4��R����)�U��Q{�#==퍜��W�M|d�^��q��Sj�'��hS�[8#��{��apz���{��3�~��}�+=VO{}�g���.�(��2�s�dݽ�Ý�=�A��fo{�-�I�dZ��n�l�R9��kS�qi�Ѡ�/��943ݨz�"��Npx˃=�|��ҷ����o��� i܄_տ���~��w��_�ڷ�Y�KBv>�UN`�; ������M�΋F��2lSUʠT�t<i�W����������y��J}�obo���B���&OY��M��mtP�7�hζ#-Y+2��G��*ݽˈ7y�=��1�D��c �ZʧuanM_ۃ�w_7�0���J�M�J�cM�3Il1H&�3��K��^C�%#%ؖ��힫6�\�� ���:��v�N*B5�f�qd���yݼ�����w	T��9�c�<v��t���9���y��#��n�����<]���Ծ���Sn�ݎ���
��Z��<��'��˚�Aݞ���1pͱ�x9f�)s)lD&�˄λa�,[(q�v��6���X�RmGSӑ�LZW�^��4����q���mٰ�퍮���sv6��O)��;J�Q����ip�^h��F�[�^uǆ�Cգ\v�q˥�v�%�t�\�s��nBg\�0��h'c��-JX�6�\t��2Rz�8��'Aw.b����s[�@`��������9)wZ��v^X�cln����y������l��� ��ܶN�R�Bt�[�\����Zb��L8�0�%[�\�a�0\��-[�e�;���E�ǥ�n���/`F���v��b�qx�u�����n:/sق㵗�θ�QFM�(�XPd���\��/�h�B�[��6x��.�z�U''^�����5|�b�.���C9>����'�Xz��/n>'���Q�͘/$&ߤ�nQ�d�2x�ni���|�S����g=��b{��(jcF6q��zTU)��)DTA'r���a�@H�4,�jG0�ίx��Z\Q2Jj!�;�K�H� �d�GO� AWv�n1@�cE�9��i���I9�Z1�[�
^(��̣��n!�[�X��\Ø���Vd&��Wn5ޥ��+��.��rw���r�#tH8���Y�x� ���U܌��o���3��m�,{�9����!$�f7��2�Hm��ڕ1��db�,�n&��H� �l	����#� G�pйRLӘ�0�px)�7�g�a� ��Wǎ��lN��գi�m����ij�f���è����nj3cżt�O\���7cr��Y\5�Z����7�n&Mh��sA�9�aK+����IV��ٲ��E]�	ly9������4���0J�.X�m��tZŅPm�b!7��Q����nm���p0�4�����ј�s���gl1����P���F�o���S*k�f�灔�jDM| �Pn�����cݏq1��Tn<W *�d���7��5�����N��.��뫥��4�TJBi�-�ڮ7��������?���O�<���\6]��¿�K9W�[��pn(�A%uwzwS�D�a����A��>��@_�׵��{�~�SPE	>�EŜ�5�gn��|qU�����nm��h�.)�0f���2�k}��o''�߾ �:�gkP��u[E�� ;*��G6�7��� ���\{��s>݉�."$폾���yu@�>5Y��#����s����n�R��T��sۚ.�BI&nUn����\�k.�qU���> ��`�@P��/���wwyh�%x��s�B=p8}�b�V +�1 ���P��]4�F�D+ ƅ�a}��O�|�T����79� W����Z,��9�Q4���6r�lZ�������I%U�|=�3��q⧽ݺ��1�V�ջ��ci�]SjuwRW���-o�B��mر��1F�&��z�5�őEY�U��'��W�ytUD��<>�o=���Fp�I��-�\�`֓���70ŭ�(*a]����>������;���s���	�ay"�������l#Q�M��n��
�pe	���y�8�~J����|qT{R�f��G�#��pV��Y�r��뉒yN��׳An� �UH�fe�Q7�/��~�>��.��L�M����Zў���ּ��t�����.i��7[f����p���I��;�mg8�%�n֍���Mv��]X�v�m�`�	g�x䞒�s�O7qá����+��Ky�-�Yy-��'e��j>Q������āMXP�(m��d#n;V�ץ�v�߀Qt����,A��j�#��(�QO����B�ˈ�9jU��y�K�A����[�ы�V�Q��*���
��{��c��*ğ�ڎ��e�8su��@���g�:"T(n!�:������ﹻё�"EABO��LN1��F]��>�QP�gI)�r囮��uF�QF:j��y�NpD�Y�ܮ��Ws������p���I����5���c�$���A��M$g���ʄf"��.���<�4�U^�ﾜٓQ�%���3t��ы��T���y�*!�6KM��DE�56�{�>=�#u����˭�����Τ}P�� QϢ�m��y����b�c�%E���8=�c2��Y5�~�ε{՗/.כ��s�ɰ�)# I"�"I"����oغ���*� G���ҕ|����ASl�&��φ���\�#���e{��Ճ.��r��B�b��2a�i��Mqv{����hpDUwK5xB��kˀ2��74 nwڗ�,DEW�f���LTx��U.l��� F(7Igy�Cm엾4�&]��z�GY�9Gko��]/�,�7�iu}�δt;� $�! wG����Tr��"��i\>�l���5�=X��peo,�)��WE�J�]0��4S��;�ݡ�=~r�+EY���j��|���8<��,& �Dz(Ah�BO��N���y�����	�8>�B�T��CM����3ѿ|+8�Ϯ_{��ޞg<�gu�=�����?a���7%NO�,�6Q}:vD'f�Wr�42��6�!�E|���2��l��r���qqG;S�mW��r���Ş9�����);h�Fǖ/n݋�n��v�7i^��&ƭ�s�b7Bc@����	ʹ���04�i��*A��Kd��s��,8�p"{���}v>��J��}���tQix�i�����ñ���s��u���[�|7g���.@,�!��U���U�(i���q��L	�!�: �-7��wp4��ޏ�R�[W�t*�Fx�g�,�m`�W�ｹ����DV���ghyB�J9ʍ�lCj�W���]��m�(��|b��~�Q�� I��l�4Z��!_4%��"�mUu�ۻ���U�5!��??�*�H�u���>�P���
��.T�E}��4rҟV��C
"�p���D��l�x� O��h�d�2o��������<��"#�i�#��.Z�=l3N�q�?����%��}1]���X�C�������;j��'lt�IS��ӞZ��Ň3&~�㗆�h�J����C�t����}?i�3n.�|��i�����jwim�<�2���%�1+{+�Gksr��3rpr����;���;'D|��ˉ��c�&|�$��'iz�Ou-b�`��,���n<�٨y4�0��t���F���yQv�Gs�{Ǽo����Ӵ�-��֕��}����Onگ��E��O�vi:oW�#^�Y�^��,��}b}3�(�y��?���I�~�������q�{C�4w�B�.*y�c����YYGa��ވ;b���G2)���9��t�q�Z�.eZv��ژ^��c�U��H���k�w�8%�ǋ%�������������	�P�mO�/~[_�4���s�\U�\%v��Nl)̖�Zb���n1��"Q�q����gw[��ȝ�v}��$i����p�D1J�!��Dr��KixTJ�{��w���A���+ʏ�`/�0�v���^��X&�.l'���ÀmKuC��-�0xp��9�����8�/6�����A���U�9����~��!��^�y�Ӗ�ss�I"V��I�}D��Z'���</�?y��ɞP�۹簏�7�tXP�3G����QI��	$�j&�B�Å��54.>�@����تŧpUdM�`!��O��U�
�Y���)��b����^S
���:;�Vq�9�{�S:�����[$Vs��G12�� �Q��#8�W��+�9��o�&����8�pY*�j�G��C�S��2��P���h���C㖹8a�e�܍ VS돴�������!�C���lc���3�(�-�s9[����;���9�u`��\5�}�.�5����43īn1M�6r����� �V�bi1U���U�^�*V��y�H�*���F��Y�����^rwiډѕ�{Evn�ۙ��Tfx������@���? H��'������;��ל$�Aq� �xb�)((D&��m�۝\� �˸���K
�ѥ6���fַ��$Jp!���yk�|�F�S}S��x$��t{�����/�3ܑq'�/1�Q����(���ܟ�Y����,�b����_�Mlɸ�<Ҍp���6%UO�2M��7�Yt���`��
z��4�V����摷��N�S���&*�.
j���غ2��u��O��5�/�w	���c����q6��Ko\�u/�宽��v.d�o\zXKs�P֭��˄6sq�;��.�.Ae6� h�����NO,��cQ��=���Ƿ��x���^���v���qa�WH�'�4k<��J����3|�^ǁ�Q#/��ζ=UNk�?}���� D�r�ſ}��l]y^ٸ�GA`�}��\֡�����Y6#˄�J}�C�}u��2�|4X����x�4�f���rH<p�I&�E�ӆ&Z���O��{��<}��F��S�λ��Z�(���P���K�vgoOWu.�����gF��S�މ/]�*{xo˾���C���@�.k��cd�͹��b�>?>����]�?�ZBSY�<�W�}�ލ�M� ^y�ȗ���Ws��#�LC�^��'���B�{���(���]Â:�x��@���N1�-��oj���Z� �v���aN{u����=�;6 yV=�'*}�A䉑�W�ϮE��V�M3*�χi4!��S[��^l�Uj8�=z������j��m}7��4�*6ѫs]�U�  �>$G�.�byE0���tVR�yg���Eؾx����p&�אی}�]�����"���+1ЛN0�i4Xn
����w�)��ыш�5~Z>r:�uj����""���}��Ӛ�:��AY"w�?훽^�.�+xJ�c�s�s�qy$ࡷLy�B̤�̸����L�CsL!Q��A���Z��k�]ݹr�s[�j�nlj�>;����<���A��\>Zǲ:�XkA�D&�@ahNT�kv4 ;k���=	�Z!B�{ɓ�C���AM����	��v��,�^�]ش}0x�aB��0g<��>�&�,�$����UZ������	���$�Q��W�Ώ��O��� �Οp�S��2�U?X�"�q��O��.��":z��o&��>����l'�o������Έxy�n&�9�Vg�V֭���Iv�٧���z�d�hK� H8	��s���r�F��-��r��0��[<)펝�.Ba��m��@�;?R�r[��1k��Qr�F�ۚ6wj�F�ݨ�sTmˮ�use`���!/%�ܳ���s6�-0Y��/g;\���6M��F�lD/�����'�q5��~�1���9�#�kd� ����4XU^�(����ķ-���S��'G��zY:a�+ r��P�Q�0�Q�K�r�}�#֑υx�i	���|~g봤�ػWa6�6��4��ߗ�ҋ�= Ln%W�|�TUg�[9��Z��r(��C.����&��e]"��KܡH��
f����	 �ܴ\�Nv+�й���b+�lTZ-r���u	�A��'�.V z̯CEBFM�9k~�r�EϹA�Q�����z$���!U�3�_z
�}����a���>13��/��"'���ێ%�<�Bjћf!���i[[,�/��}������KD��y�>KbJ�����^N0�J���˦�M\nFlA��Q���"�X�h S�Q�fi���Q��I۾5L����-}#�;��N��ѵ�᫛t�#1����iݎ���\���bJ���5�ߴ\߶\�Nn����S^�z�E\��~Z�s@�g�h6a]�G~5�O�-J��័���M�jh8#��a-i�p붸�I� �U�,�%��L� ��x-q
��D��Н��Q��|~���H1���}�ՠ��y�O�k���E�U���a��l�ҾW��b����+��⪻��5WH����1���E]�)��,�k5A�n��ܰQ���m��nW*�ʰ�HDFB��]�y�xpԼ��4$� ��0��PF��̈>&_���M��r���.���!6M)��Ϲ*�n��}�qܑ�B8(��#"�ɏ��a8��gr�#���>�Q[��[�p|a�^�;!�T$g y���J����H�$��yDDU�#�L�Z������y���������a	>rI$�`( E������?˟�W]]�Mj�[�Zi����0Q-���Y@BDAR@	W�EUZ�(���X�+k�ڹ�Tck�Z�<*"64TkX�5F�U���V ���5�Ebū"��5X�k�+6�mEE�m�mQlj����F�cm�+�4cU@m���ыcQ�m6-DQ�h1�j-�b��6����h�ƍ�(�	�j0����,k���Q�X*#�cF#*�TZ�m��ƨ�E�(,[F-A�ڌU���Q��Q�[�5�ڋh�V�hڊ�DU�¶�b��kkM�RX(#�T@�(@�S���m�Q�����Z�F�Ub�\�[l[kEUogM���ŭW5���a�@!$Q�R�"�"�����Ŵm�.[Q��Vf����i��u��Ƶ"(�EPj�FP���@A�U7�"� ���Ip@j*�lUDȤ�	pU;�|7����T#���?dTEU�IFu�(����?������﯏���?����O��~���������X}D;���۟�����[g�����p��~?���A��(����?��u��Q ?$���<~?���_������P@����?�����?��O��h~��
�ߟ�E�}?�R��O�S�Q >�>T����~�'�~���#��?@��q4�j��i6?���E��	T��o�n���~IG��@/�s�1�R#"1D�6��֖Z���SkM�����A"��$X��M�4���֖ͭ*�	"��$T�$D�$mim�fڔ�ٖ�Ymb�B(�"�B(��Z[R�����ږ��b�"D��$D�E@�Q�E��X!�$@(�A�AQ�$X�DP�$@H
@A�$@H�AF(�  )�E)�b�`� b��D�E
DH�A�EH
@X"@X�EF � "�*`�E�$T�5��������Z[SkD(�D�$Eb��ER�Q�$Qb� (�Q 	! �P�T��QH�D"� �$PF��E"	�T �(�Q )(�@`�Q�Q�$E"��EB@"AH�@�@#"��$F(���֔�����kJ�eJ���Z�m��ڍ�ZikJmi���j-i�m4��6�٭���i���eKe-���ښj�-R������,�4�6kM�-�6�6�*R�KS6�f���fm���+)e,�M�YIE)��e2��JiJ��*S)�%6RԥYMf��-J[L�SiM)�������R�fS)e)JRSJl��̥)M)Je4���QV(�Eh�m�2�շ-�mXֶ6�km��SKR�ie��ړmL�R�$*V �(��$��Vk�@�Z|��F���~�ׯ�����A{�4"ڨ��b_�>G���7�����}����������:�/c>(_�� A�� ��R�-=�~�A���0>��o�O��>=|���߸t������xHC��'?�:�ߏ�'a�Q =��+~!�����������9�����������Q ?0��_�i������h8�_�S��x������(T ֏�=i��B� A���������@[>V��e"��+@��%��̸;Q %ſ����}I�	�_�D �Ck�������U�R�����C�����3У�8/������{��ŏ��>���?�~���A 	��a ���?�D ��B/ۡ���t?zv��C��#���~!uiD�q�����>߿�/�����B��������(� >A�?��Q�����O��m~�:=��HD�I�~��@����P��Y��b� ����}_!��b/�OSo��?j|OA ��8�"����K����T������߅��A(0_��|�_��ܑN$Vŀ