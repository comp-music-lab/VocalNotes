BZh91AY&SY���
�_�py����������aA?4 @   4        ��    ��   }  h@�[4  
 
�� h >J �U  ��@P�P@QB�� &{�   /z�>�&�Kc�Ӿ�Ӡ!�wE��{��mC+U��w��
 @ s��wS��@uu�W�OYc�w��cov�L�y=������u�m�8���5�Ar�֝ϊ��J�   (;�(K�"��l�����zw�y��׷t�!�y�o;��z�ս��0^�G�oz]N�t�<=]�ݱVv��(��o������m�Θj�ݥdn^�;�w=�G�=��w�9��s�9h�{ۯGfئe�>JQo�  �
�
^��{�̐m�����3�n	Z-�]�M4��<�:]�1Xg�T@��Q���r�w)v$hv��2�ø#ttu��a��	r�Ԅ�W�� ���{û�������^p{�X���7�u�{��	YwnE��z�*
-�����Vأv$��@��ѻ �N���   P w��̞أA���9a�2:4�����v2B������:������E�jՆ�`@ݷb����]��                 Sɠ)J�i�a1@ɀ� �E?R�SFL���2` M10��USCA&`L �0D�*�BQ    1   =	�*��2b� L��T# S������b�S�&��=G��G�}_?�}�vk��~ "(����

�dT~� T���@2#?��_��@������4J�r "�N$��|q�- �'?�	� Q@8�/S�C럷���� �����<�?����b�mc�����|[�����@ӑ�&�)���r0?�F��j��},�v!��M�g�c���2��S�+���"�(�l[����}I� �nr<�x��97��5�����H]�
h�mvͫS-rd��f�sN\r�΢�G�(��@�P����w���F^���VM1��)G��t�c1
FϦ��ρxw��̍T�M�N�{.��D)�p�p���݄A�vr�.�4�{׸P���ئf�o����=8]ݼ�NCn�4����x�1;vD*��	؀xE�����dt��sx���݀��W.��5c �Y�^i=OK�N�}���u<�V(�^�8�b�[�va����Q��$��E#/T�.�Njӳ�`]
䣗V�����IMl%�cBҴ��Y��)'���2�5拚h�i�Oq��a|y�s7v�*r�EYײ���)������;Mm��E�c�ҧ.���p�аN��+�T�a���[�t���P�V�X���	N�#�^O!�؈�;����T����砅Oݴ���<R<)���>��G[%�$k��߇P��T�Rjgo)�p�9Y�)�e7��pѠ�\�s���]r�A��ۛ�����4�^��Ň�]N����e �0�x����kpI�/%���$��ɚHY�a�>@'T�7�]{��.+�$'�6�7/"�xH��h锭��A��ӂ�w(a�v�T��˻��3�@�)�og��O����݁�c��#[����v�2��\��s&־��������j��iU� ����u�+ӡ�^�l�����`�_�M������XaE�6$x��;����_��:�h@�P�f�\4i��T�4�^Mգ�Wqs�l�q�Ank�'Ut�i��{+ǚ!0���c40"�����+⸎S�c�'+�]ݗ�\ԍ�D�PWou;����n�2m�/ݜ��63+�L�З�t�� �ig8�E��ߘ��K��Zj��J燂1�ظ����yv|w��k��-fH8r.5�0u���R/9���	��N�T��w��^Sm�I�a�C��� b�u(�q���״(C��QG;����˛Wpn�{prs!|�z�+�A����L������0����A����B���Psps-;8�,�"��2�f�R�s@]�d���{�vaU����z�8X4j���dM�����X�Y"��a��$�%#�����05l 0N�
E.4�L��Êvl��OJ���.��ܸ_=&뙻��Jq	�����e �b��A�;���w�v����K����&�w���A-��ײ-�Ĉ2�E��BVp0���%��*��XjhJ���sMǚn�y�#{�p1n3�%��M<���A4�-�+f	�����נ}T��H����)���^�u4!��ɸv\��d/\ ��@#(�^���蛓�z8�X���q՝���v뚥��v����y�
�H�Ď�9-/g3�H�p�QKNi�-"�.ٝ����n�y�m��q�G��ֳ��f���gs��0x���z�t=u'�f��[�G�uqL���7���f�{&�I�JF�rTf'�5�;���N�j�ɲ��wjfG���������ns]˴l�۶^!@���Aņ��Zu�:W��W����rwe��<Z]��@�;�����*!R�)
�@�ߧ=R��t�=I���,��8�q>��Gb0����nn�M3� 9`�2�����gp�7�O� ����8���r2��T�<Kzvm��q`���qt,7�sz��Ԁ\��sn���w�jn��ܺ�\�j� ��<����Q}r���foփWW�Q�bA��.Q���ieǴ7�N7�Ͱk�ɢ�'e�loJ��s �8�.��ŹQ԰���؞ۤ�!i���]������i����pMrs�{��Ժ�tL`�4�1*l�׵^���������zL=��r�$���Fq�>�P��m��g�ٯ��b��#�/i�����ҟc�Q\Dt��L:.f�������)�&*ZѮ[@N1�7{zw{�]�ڷ����B�	��F!� �`f�8����f�#-����VН�l�K� �6�Н<�w�-�ygJ˒1&b}��F"(��N��5�d9v�hLә�ة��yCy�nM��D��NW��jJ6�_vv�R��6��;��znG_Q;P�h�ֽ��2��r�bᡮ���k�����<�I�	S�;�G!΁=Љ���,�4��0��7�7@�k_Qf�;�q+�(g�9n,��[�i;����0�q��+�O坷$��Lk�M0���+E,�� ��H�qC�u�v�5��GB�T\�D�rf��D����gp���5��{x����]��0�IIm��vN�r]���{�aF�ӛWe8�0/j��8���zDt�{7/'c��*��ưb�Nc\��%�`��b�b�;{v��qly�KiOw
@G�0־Z�&�n��ޭhn����䃢�܋-�ݓ��	�Oޜ�t�7���6j̃3�X��ݓ�igo��h�>��'�Vyn��v��C����4��� ����r�w0Q��Z�v��;p��MSX��K�%;KR��Ü]'-YUQu�g�G6�Ж&:GQ�m��,<_NPwʄ�m
�ޗ���Š]��!�%��ۦ%�#-�`�DcxT�9a:�o0�e�f9q�"��&�t��c'���36<=vR���j���:'n�u�.L�i4GqrkE�nv�ۭh(5>O��� �f��M݂������=��Q�.yA�(F�P��4�����"7�dZ��a{�)�:�\���n^�^��Xٙ�sm��o�q};r�5Z�d����Cum#�9e�Z0u��[r��]w�K�iޭ*9(��Mm�+�%]��v�ܜT�E��vI�n�ڪ�A��������6:���+��K�j�F�ݛ6a��G<\:Β$P���*�}4!�{�\�lT[EA�3����7f,=g�dk�1ÕD7��xD�\HrYOM{�m}�J�Wvo�f�e뻵��M3 owpv0 ͔gi��鮐�KV��h��ٛf�>d̨^�w8�4v���[��7�����k)�iF-BLRn�ݶQϏ]���&@���r��{N���B���ܸ��_s��D	��d��S���eN���ڎ2,y5ν�Ĩ�׺����ܰk�,�?n'{��m[�V��u�7g=Q��:;�8�=]��B���5�Œ����6�@�2-]6�ۃ]E��:]C��'�n�BY
V�&@���ۑ3�C���]�5��Ax�����Y�t�]��'\�J�٪m�t/�D�h��J9	�GӜ�}�:��be���� 3Ӯ7�[�Z鍻Gu�վ�]��Y�p�7��{:ps��=��N���n�{w,;��dH�:�"�Y�.ḝ��7*sw؅:�Ĭ@&T�^B��ӂ1�S0rrV�80�ˌ�U��c�k<S��G�Z+�U�#M�(��C;��)�{���C�u|i�_PL�����H1�]lEPLT$���`I�P����-ʟ}Q IL�.��v�1�i{1����'p� �7%��{]{�V,���5h�2M���\�gW�Y闸gr�ý�����t�?{s�k[E��1qX�g��V�^�$f{!3Y1����U����Q_���W�嗡�N�G���}]{��Ó�>��}j~�9WK����Zs(�k����"Gcp��Wln�뇶��������uXS�^q�k�=&ںh�bmKv��\��5���r�%��������z+���ֺ.M����s̉�r�q��������!+���y�خz�uR�ܵ�t=��`���6���1�n�7`����6~5s�ە�r���=;:�|V�vA�7/��c����ݸ,�:3�m�c�H[�`j�01`#N�n{p2۞���p���=h^�Mα����'1X^�&(L��Y9.7>/E���ثaypܽ�����hmQ�d��4n4��uq1�d��x�&ꞷ"H�*Y�P��=��$�m��9M���]clrtnn��K۱sp��PI��]��u��+,��ǫM#)���ҁ�:�GsƻGۛ���<a�"Hĳ5J\�dv�.w:�Cv��<�!P���i��m+h��ȫ+j�\]UUt���i���X�oKs�5�i�n�j��=�svYs學[QA+���Y}�Z���Rsykp��s�vu�'^oW^�{t���e;jk�v�1���l���t�#v�ۧYԻ��0��غ�o+ӎ5��J�g5�/+c���[���8��Nл[�,���v#d����p�S1��җ�nx���#��$�!݋��8�[�� �!N���`u�ںpKΟ4�	�wa���쭥��3��n����[۰������9s�<��6��ֱ>�6��ne^�!类p+��p�	�Ω�rlsm��K���%�n+��'��tv5����ۅ��Z�I�s&��غm�2�T�]�������1���GG�J�C�&��2�"�' Vj&"��^wVN�D9,e��l{h�n@9��<���[�2��<%�l�p;q�k�s��z;��I��:�v(�/]�0����N��<��u��R���a��bxW��8}�d�v7a�C�6l`�x+���9�`�`��V7=�.�.�x⧢!��U�D�P5M�z��	*���ƴpOclu"�]q3)Y���gm<�<��Aº2)t�O��+�����s7eG[A��/]���6��:��WV5�<�S�k8j-c(�x�gk,�/={�.�\��͓Gn�z�����e�"�r0B%��4�T�,����1��6��-Ŕٞ�R\c�[.��7n����ࠎNؔ;c]v���q
��z��Y�ϥ:6��ܞS�}_�?9��>���\1�d��Y&.��h���vщ�j{���䵍Y��c��Q�4�#m�(��Z��w4�M���O]����E��0Q��u��g�^;��I�{�u�Z�n:��+L���Q��ֵ���1��������)0c�`7�-�f��r� �Z���ۭ��Y��wk`�۱����䌠�� �D+'H�j0aا�^��s���/��LqY�[;ƣmx��u�6K�X<�f�H�ǟ��/k��_
���m�drj�\�c����Iɾr�'
�Қ�n�uLr��p�m���F���B1v{��Y]��׷]��\�pݶ]��gt���N禛��A �86����n�qYv�R���9[A���wA�۱q�p�#�O]�X�"�Z�;���^�Z�gԼ�$�Q��*vy{q7<�u�q�pL\a���ɪݎf�G-�	Ӳ=ό�vu��n�rG���Hۭ�"F�v�uH%g���'��]��n1�L�M6�76׸��u����6T�Q����s��Bt?����?Hq�˅�+��ia�ta�oLd�Z�&ю�f�S����v�Q���V���UBr�bn���h�&�����/�1�&�rW=lr�s�獋2m�C}[��\��{<��i�4�˥��u�b��q�8/9ܚ��=;���vve`�5�Q��&)��<�Y�N!.�Y1�A`�k�ѫ�8����胴�q� n���ֺ֝��nϮ�{n�Ҧm��yв��v�F�h��u�s���>���/��n�0���[p�^��J�%wt:�2��d��T� ���8�p�������|��g@�'7@ˬ[wR��`+<,q]�e���F�ڠ�F��ʩ�q��O��qC����m�����؀S���v�	��S)J��ji:�"HƓ|��/o���=`��)���ۍ��N�@q\���F�R�e �DSې9��)��/=���Jjў��%����]�i6��t�nkr,\v ����<ݓ\� �y�;m��>S����#q��n��u��]��,�5-�*�ADK�1�J�J��d-pnT$��*�\�s�7m�\���s�.�sy����0��<���n_a�a�W����=q�qnw����)خMiw�!sp��y�KYD뉎�h��E��;\���nq��]�W� m���VtI��i�qE��V|x0��p������!��;ү ���5�ݮ�6焻��>b����૦��\@��eb6ܶL3�8��y9�v��Ǉ�ɭ�;7�Oc��1���m��WA����	��̠nM�-��0e��~B�pn��Әc��ܼ\��ss�q�]�lq��鳋�1"�Ƴ��7j�u��_.�]�4v��-�!��q���lGa�Ѳt����Ή���Sl���n-Ϸ��
6�>���ۉ��;��,�s�b�f�Qd�i��t�N����Wl�Yuu)!z�uf�J�q��ޚ�݆h˺�����î\�=��nz1����hF!��������Q����g=	�mN9�n�X���FmsCY���v��ۇet��s�AZ8�t�^�o�\ax\�MպL�����Oe쾝Ra��j>[�'�PDP��"�Î.v"h�e��?����_��_����>���8���4ҿ�5�_ܵ��d����z�������+v������m�f�v�\�Ӱ����)�q�w[�k3��vG�:�ճʷ��� �ئs��*^̡w]��-Y���!f/+4�����'��z{%UL���a+����Wb�}��:��G ���STm!��s����w�H��y���'d0�	�z�U	�0{&��t��*���]�s�~�����	WY�]��.�FSR(T�m�%���A��;�2�#ܽd�7��j�ݓ|b臱@�����o.^i�V�J��tC:ws8��|�:�C���[�/;|`��ދx�D��Ӽ��N�m]����O�m�{������$�Pq����#�z��s޵9���9��[iz>=K�03��c������{&�c�� X��~Z��t��[E��/w{5�cJ[��>��>�)��w�%�`F�.A潸d8�5��u��M�	{��Rs�.jŔn�_r~x�d�{��+���w_q	��ڧ�O╇/:u�i}�=��ܱM��܌j[�
ۈ-����5���/-�%����bm�����ݒ��X�i��ٽ<��f�cte�B��n��ǛRBgڼ�!��H�>�����ܘL���ݲP���z����j�G�.GT>�Y����&�����լ{ũ4�v�x�_n��c��~$^��)����&����c��k*�Ј����ے�#)y�� ��)]ں���JH"s^�a����9���{0��Mwl� �Z5����zxN��M79\��H��O-��H�w2������������o�p�6d���<���h�Z3��;�u0=��s��B�5*��s[������5Yb�WrDQ��'�Ϩ�3�S��yM)��7�/��iΝ;��bJ[v8���ʷD<��Iy�~���WύX��/Fm�������f��t�M���|�-��&���k��!��0;�m'
ȴ��r�=�^(R�>c��&>�麌]��u��͸ﯔ���VȎo�����ı󯷧�Om�"װ���<������}��bz�͆6F%�ҹ�8O<|c��;W���gv����3�p�)����B�tsk�7|�{����c�ov� �>�]X�,�g�Po�:s�W� b�'A��u�t�?]��m�~������������yM&�wS�or,��.�
K��n���:�<�pC����}x�kD4�/9sGv>a�Ny�t�y�z;�|�pe��4��W��Υ.��Hf�kw��ռ.U����qk���ǃ���Z�U��R!q������8�xi铄��evCท#f �giL��4�p�1�j�uʌ�a^!9b6��Ë</���v������b��v,'�
���Q2f #�ӻ=�o[5H@W��y�i��|�����n$��T�t{k���Q���N��D}MT�3�HW.�^y�94�+��;��+��1�0���n�j����]��� #�\+��
ް���N�H�H�u�s��v��A�f�b��e�����!���we'y=�v�#�<Q$���-Ԧ����V�g1�Lc��fyUi�m�{�y���[쾀���[�tj�O��>@��&����O�swS�S��juK|�HU	ou��Jw�3����\[������-�1���R|�9�`4r��<�|������|w�J��~An��y>�t�S�G�p�͆�DT���zi�8M2J�L������{u�΢#�Z�Jx�W��K�8�����i3�����[�hW��zps/�f�޼�|;<Avz�;�_4.y/���ɳ=�!_7f�1�4�<c}EBwhvOZ���w��}��W�f� �Y�m�}O����n�eW���_ܸh�!��g������;g���8�B�2�B��z���#�:�C��{~R5̼�n!�,�IU�ףK��#
����bf�jbq�l��c=��Vm���=;]��==;�|�[=	~��U��N=����.nO|���:��x�	,}l3'g
7�;+��d�wm������|�/��wˮV!��yvH�l�)��o���g�\+�)�׋=޽s�nw�ؼ]:>�����<��佛�J�s��K��8�{xN�Ș�ѵ�e[u���V�H�v��z�(�y�?#�h�St���K�c��ߪ��Cz��7�ü��7��@pU�g�<�4�<|g_p�.�p>1{{Ze^�g��r5���<O��v<�d3v'&�H=�����a��@�B7vNw�����Q�-%LY}L���p��4�w
��[�yIꋠ]�����4�����Zģ|��f���g��
���L�W,;�F�p��n?7��.x�)���y���>�μ>���{�g��$���{�)$���o��l-�P�F �m�������9s2w�g�=}s�*$\}����)�q���y�����y�j�OS�u.}�ci`����C���{I$�c�����V6xc������Z��g��0��W���v��:�oˀ�7�����X�VP�[9��u������-����y���s|�;�)�}��鞆�$cO�8�O-]�����:z�6xUT��Y;پ���W.������ţ�{���Mؒ��?0MK����Sy�X�1{8=�0�F[�!��y��6ZgI-K��F���.F�ެ��$QD>(Y��.&���;��gj�p7�����g���0�w>���t�l�\�,�L:Ҷ8k���|��0v3�ݻ��RC.�<��}����y�B����+r����S�4����+b����	�N��u,�X�V��o���ټͻfօp��Ku�:Ë�������]���T��?l�=�;'�/{*����xqG����&vn���8��(C�ť��vx�{Er{�y0������I�E�Vnj�J`	ʭ��g���Lf� g!.$�whM,k`�=���{H�����,��ȽL��;�=�V��w$�M�8&�,���6���S�s�e�}�gєr�wZ�QC}U�#�ݺ����� ک�ܘ���w�gm���=ʹy��˷�v�Pc.��N�G�/�2gs{g��D�<<���U�~�Rz��Ff��z��N�r�H�����y ��۸Щًn!�e��"������1zi�S'wa�.R���-�[t�7�@�3*X�����ͭ�+mȢ׍MffS����;��M��	k=3�;W(x��}{'�o���yaW��_�>���A�@�^n�nd5�*v�ˬz�t��Y�ٳ���>[�cp�ҝ�Җ�-5��ޅ7^J7F����]��⥟b�=?PJ[����j����3-b@4L$�=n{�<�FD�=��p�{�h���d�ǔ�6��!lc�"A�Zx��L����9j�Ͻp�:3��]�7�ͯ=�q<�4e����|�8�LT��h�<, g�v���~z�9�b��_w��/TwӃ��:���@"�Btxﶿ-k�w�����0懋�b���=���ڼ`�K>�-֯�s{���p�� ��\���Az��5�?u~��s<v왻�<:�ڻ���yb��w���\wS�:�$�^��`Gg���<I9�CL�CA]�{t̫&��gx�AQd�{�[Vj;�競H;���{
���)?2Y�iM��-������EZ=�w��b��nw��F�1�������l����#�	{.um���/��F2�BzbT��i�{��,�4'�S��׹^մ]j�QP�v�Q��%�Ho3.�����h��s�'��|��G/����߻=��{�i���{�z�=c�������} P%��=~���>�@�����kX�8,}n,d����j�M�Q�+	]�%�]�&N�6�8˷s��.t�tF�]	*���<��6���N��ո�=%�tZ{)�0��7N�i�2�91�-uڞxIz�=�W��(g��ٸȔ��͢��,n�F3�ӹ;x��C��q�<s���n�m��Bts؉_Vx��z�9�C��׵�������F�x����z��1nN��^�tVyv �k�V�垸�x�����r+�n<.��<��>z��m�ui󞮝	�1q�����c�s��v�I�:SZL�m�1�Yh�#6��6Kgm��Y�s��&xwD�)�����[a1��x���=r=����h�+�gu�X�qˎ��8�q�&x#�ɭ��n�'�y�t{�NN���f�^\�Ӯ�Ο\ݷF+a��n@���v��v�����q2+ѳC���\`�qwj�9�uǃ�i���y���ld�]k��f��9`f�<%r���ۅ8.v�����m��v��]ĻvY��+ͷ/C���h�ہ�u�]��v'n˨gP��l�fi0�;fΘ'��m�<��Tuj���{3_������$%���%h�Z�x]iW��輕��h�yj2j܍W�͢S���õ��ݲ�J
F�%�I�Dcmn�`;��H�ti��Wp�c��Y��A�p��څ��S�﵎��"��I�S ����a����@u{; 0�,�����*p�JRb �ma�'ӓj�|��f+���05��gwt:sYtcT#hቂ�=Ҫ�	Y@oNԺE;5*9�ܯ9Y������Wv����ǻ���6�C��W���ڜɒ<�w������[��a���y��q^
�i��_���&.�N�z��H�h�[wa���m�=�����+���Q˝ő�o�\[����\��o�0��%a�t��]BЊ�qM�qXAuV���1m�*Ř/��)��ktՅ���E����/=,:�H�S��y�%ck�cQ⤄`8�����h�`�����O;�7��I�k�Ӂ�ᵭld�q�t�Μ���=ֶ9�u������te1h��o=���������:k�݈������X|��}ס�xd�5>D�$�u'�!��j6&�Hr�(��DwmQ�C;���؞�7ѬB	���8 k*�ڃb��C���#3����������3��@2HLBP' ٓ$���B-鎽��D?@N�e|'2��cW��ėrp;|��Z�r�`� ����c�t��r�D�g=�[�i�*�3�}�p��҉�̆�P�bM�7w:,�܋�9}@'Eu$u��u��sr�w�q�ˉL�[��q��d�qy��j$2�j�z���V*A��H�^j�� ��O1qlx��ڋH͝�l� o�0H}��ը�	��(���M�����b�7c����M���/�z���8q%_~Z��UTq2彎۸�;z�\8�����s0��3�%VdM�-�5���G&��$����b�7[�"E�v��DC��*�T�7Q�#��j�N�2}�C����0�u���%��nz��C��A|(�>��,�$� �y\�2�G$^k2��z-�u�q�A�2_�}�k4ov��f��� ��%��T&��	�e��	���2������k(d`( ه�����ɸM�{��(���5N�:�����N�$#�ʔ����
M�Ͼ�񩹮��z�!SZ1C0� ���RꞞ0�nt�Gs��f�����<�&����fǯѯ�Q��f�S�VWu}����A�#�o���v_6�u��e�2'�����,b
2sLJLA$i��&���Q�T�؊0��F�H� Q�<���9|$��(w�"�tfV-i��U~=��\vպq��ێ&}NN{^30D18v�lC�a�UkG��Ȥ��\"�mƗ� ���fM�����W��d��yf�ehBj�3�aF��qt�z��G��vnHzoh��P��kg�{�[k�8�ճ�z�V��������(׮���\�[ֽ�;���7D9��.��^
%0�q�dxup�c�ã�ZR�]��[�3�����+�;���*��{4�Ǒ,��w(E�X�3qm�Qx���[�
'e����B
��@ �nu�C�v���<�G�� �R�ϯ�+F���v���7L�rf��Z����O w���-��8����]��'V{ˉ��Ё߾׭pF�I��>[�`Ä����;�V{\(���{&5rhd(�i����Ʃv�J�n�Y��	�Ew�Dqp��mtSE��
jEy����#�{�]�v��^kW�(��� 녕����ȩJ;)+	j��h�U����^��b�=4�� ���ɡ����
sF񑴺:#K�q��V%E�
�@ꎪ�#&�]�$���:��r���
Fj�w�؜�Di �wS���ũ���
/ A����{�@l�F_tA��g���ljE��`�v<.;�Au9+�ٓ����~��p�m1��['������:�ڢT�@�c9s�Y�}�����۰o��T�[ݔ;��q�����a�	R�f0輐ڨ�ad_��u�@��%3��"N�\G�GL��I���:{#iLN�=;72]�����;41��T�Ԉg�뿅Q��I9껎9����&
$�P!>� |�ԇXQ�)?}���+�"���e	=��ash�(�]�yg�H"�-�!9�aUi��r��sťz��!��}{���!C
N�E�0�\h �MզЈm6�w�4x�f�q�W��]�/݈3`h�{�<�+B���tY�BB�mq�μ�X%��<��r�N���uF\3N.�(�+o7�����u=N?���'7K������Ƃ�|!X�Y�-p������7$xq����6\�䮵�6��v&

�E�#��<��,�Os���A�bI�XV���O�
���-My'VO������\Vf�1g�[9P �����p�01
elqmo�xSE�������9��>0'a����w��ն�͌��,�q;�=�g�*DLs�������,n�J�P�i&1�p�Mm�m������c��o"��-6����u+]RJ���h�=)6��s�w�]b�y�]K��e��ӽa��UV�؎#��,x�O����gz2`B�H8��S� |���EN=��Z)�}wJ�f�N!G�@��=^�K^�sg>#��:/����w	��$Zߏ�f��=~���S�E�P�[�'�;=HD������0�%��;�a�����s����"��ą���n�10���4^�]�EV�N���vvs�S�#-LN�R�!bpV���^�<:`J�DF������(~P&�xs�9��w��8�����"J�B��s!�wT3ܐ��je��Z*�}��WoW�;}yz�b�ר�G�!f<���&֬ �X�[@v|��'ï֤�i���,���S��q	���	�/�y����"�h���=0����Đc���b�R7c�"9��	�R��)TQ0\J�'�B�:��H�>H{)L�����|0��H�z{��y�VI�)��V����8�����@�~��郘`ď��G���Dc��`���^�^*l��E�lL�)��5�6G�7u����)�n��*�]K�4gn���S��n�pWb<������Dֆw��f�Ln[��{�QA��v�Y>s��N����A�B�f�V��Ŗ���*��LiˇV�f��*�a8��N�Xgk�wY*����ݍ�%
ִ8�è=�s�\b�����Dl!%�;&�Da�IB�6���ݚ����l;��Lם7(���v���5���S{��bܩ���r��S;�p>�U��.�w����W�,.ћ�b�'zG.���0J�1��Ӕ�`�M��Ap��{��Ѭw\25�Q�����GX���^N�P��M�E�ʌ.D���דb�D�0Q�OP׺�J����t���b���\�#dr�7a`�Y4a*���Ȼ�����5���f�6��
�����՚�	DԳ�{=�Y�kc�7P��8��͆�{ �is��ì� �K\�����=��b"�p������kBb��t+�:����z��nOs���Qc�����Rp��s�$;;�M�p]~��uɹ�x����:x,�`8Y˼�>���ݐp���l�}��?�ъ*%�^��,�>�.���M�!�e�<��/0'��E�_zamjA,z�OS�Z�6g;��idmm�)e^Q���9y"�^�D�oX2�Ρ቎.9#������������]vg�17�{�7DO���e٫��=��s�k�Ve�d�&�^Ȼ����lc;�b>���fm�h��ž&��.�ݺ=;��i�..��}G|U5���;[� 
�����()��2"4�$s�&�"�9�W}dȗ\s��Ůq�!�ϝ��X��0� a���&���^��-X�c8S�0�bt��ٔht�2<Q��ZO��^��~e@.*Wn5�X��u�K�wzz�v��z�%�j��vs��kk>�9����ӗ'�;q�9 ��L.`.8��~fV�\I�=��� �W6n��_;�f��L ��̨��3!�w��l��Գ�h�a�N�S�z���$��~�CcN}��۞��2O&��9��]�G^�t�b�������%��RB�T�-")5D�qD�RÑff|����ul^%{�&F����XM�cδ%8��6ur8(UlJ�0m�m����&6��OsEr�Ăbo;����e9���;�&P)�ty�d�α����(q�<�A��r�ˈ�`�G]��:]� �W�u�2zgь�[8Ԁy��8є^Ǵ��G�{Ȏ�]�X�� �T5 ���`�L���kx�@�N���9��뮷�Jr���Щ�=KĞb�Z�I�������LY�8��{��pz���y��5*yPI&&��Ō�:.{��X�y�Gة�}������{n���+3�@&������a���V�Qdx\�8��8�p�{(��"*k���l�L�:^4H���kq���0��\={�C�w3ܮ�\-�6�˜����5v��A���G]ƣ�g�n���8���=�����v��鑆F>��tT��b׫uJ��q��F�yMs�=��p��}^�U�Ĉ��pցbmq�.}��R�o��a��}eK�}Ǚ���JM[y��3��bYZ�ģY~�f9_<�fz�wɞ�\c8��gb��&$�{��.���P��5��x,K � ;�?{תo��#��.���ca��� ����x� 1��M�qg��9ߡ(�B��L��d GP"e���dA_� oB`��ԧ���g��=����z%�ߟ��
Z;��B��H�����-�\���{^fk1ע"��*�\7:c޲��^*~���4P2�4�!)�A�D��0Wz�-�Cyo�?�C�L@���e;�r���\�GG��Ğ��t9��9�A�=_p�k
Q�8C2y��g�6h�s�:GA�����xG;�.��#�}ޙ��Z������a�\�m#�\Hk6�o�������>��m�&���v��tIJ(
�dz�]�����������>11%�pk��G.i���8���kGs�5�a3�0�9	�=�X0V��p������$�i�DgG�G��I8�&���U�Moa����g�9��UV�O+���j��/�Ԩ���b�X��Ui��'$Ȁ����{�X���`L����˩K�2�|��2�VS%��|�ȳ�LZ�Ěy��|�!�# �$k�~����ː�.�'r�3�f2��oI��x��7�f-3Lf{݊���/]�����Ŝ�ʗg%ڸ!w=<�g����Ү��
�}�����?=�^E���q-�ŔS��h����Ecc��s:�)�������&�p�9чP�3=�x��DL�c��}	�����g�!�I>q�/3"̙g݂��y9˙^g�����7��^�`� K��2���~|���c�}$H�W��ac+��V�4V|ܼ}9���J��4TϔO���z���i:�L7�!i�(��8�p4���i�<ض?�X%�A$���M���78$����˙�3�I��<�b�S�|�L�$�<��g���}��{��T2l���g�eV�7鷽�]��4�]ۧ��u�r��I�fs�x�:=^�9��.f�����s�=��詝1zu��Y�Y����.�h�Z��雎���Ė�;쳊�s���L�}����N#3���t���8�F:�)�jw'��ɹܙ�������2s��D�Ƨ�8���g��u�2�����Zλ3O�~�L��ދ� ��q++��8�]g1����b��h���/�డj�k�/ri�G�=�Գ�L�Y]���}��v��#d�73Fȉ{gy �� \��8ˮ��&Byl��unx���pa���p��c�b���Ô�Z����]m۰��1㧠7��s��0v��YT�wEhx��U��[��]�ŻY�JYU�J�HK\�zh�3 �b0B��GLl�b���`�`(e�����*p�q�q���/�������ɜ�A��R����]�01b��Rୋ���3P�c�{4����I1$��1��زE��<�����[�E�6��e�ۃ�����6%sߺR����%,` 1s��<�ݒ��q&:�U�u�S1�����)|�ܜN�9�VCP��Gq�u��Y���]�e�("��w�]O^���Ƹ�:�t81H�Ïs�~�g(!C�i�@�=��1G�W����ݐԆ 랻�`q#���X<�Υ��u֝�RR�BжH�Tp�n 77nz�	�wGd�^k�k3�u��4�{�������C�6�.��Ŧ��J{޻Ҳ�
��i(���S�s�[U����#���&���o��
�z�2w$OL^�) 9(<XD��9;s=��Qx\�(�1N�[�@�{����F fD(�*<Y#U<N6��'�z㭎��.��̦��{�I8�����k8����q�̆�S�z�}Z8�.���uu��ݏ<���Y�('����nڗEL�ї���fG��p�{�dq=ޥs>�%��>~#�m͆�h��u�rn{S!�H����d�sמ�����!���y�?7,u7i$��9�%��3r����-��p X<�r���78%��Fx�?v�%�/߷¯ٜ3�Ȁ��~-�k����,���Av~��ٝf3^o&�Rg�z�gq9���e;\��O��׆#B!2�D��f��~5)^'�q�"m���ϖ��ꐻ�O(�%n��{�r?}��Yί:�b�g�3)��𙕵��yLt�ipKu�e�m��֊�y�s?�7��Z-2��4P�1�爉�m�_���_�}��#�:�2	��Ţ�h��Bhi=�����=<�{�g6�a�3=���v~ī�B��rlD�Q%��ۚ,o=��>�ZF�
Ё�F
�:IXq�ITM��9tSD@���g�|��u<s�s�s`�b������7T������Wޓ�"zEO��a����|��8(d�\X�L�vf�}�M&fp�b��W�V�78f�����b��v��ą \1����a<"�Q%�;��-��nrб5�ǽ� jq�)���=��	>����D=>��1�WM�oA���� �BH5�`!&A4u�箼9z�ѣ��ј�&'sF'���
c��G��QN��b�J����BA��N�Uc͵���Gev�YE�!��ٳ��A� �,~ؖ�4P��qc2��_[��V:#]�WF:��M҅�������\MێBj^
��>k̛�p�Ø\{����Q9�1r}3(�}_�H���Ny�ߖ-bJ���V1i�O��-�^��)�	'����96S��w�31K&H��8�0���EI�wwb'��¹m|"�,�,=�1pT�{|"�4Y�򘯘�Y�ڗ�A?WQ��Y�ca�fy��vMN���NY`.�ɔY�}k���E��,��'���:#��٬mXT�5tb䯓tki웻�� ���/(�V�\�j.kZԬ���{l���^�4�\qd���~Kv�R��چ)��X�[^�V�jOrS�J_��@{�A���n���=�(Ί�ٸ� \Ny��T��y4H���dZ���\�k���|moy� ���ؾ�z�{n�8�j�8*0�"�QUuM\+OqU=�B�_mx���r�NҊ���$R�r�h~�\'���1x� ��~G��������Iq귔���YSS��2�DwB��l�s=R(����s�.h�]e���Yٌ�`2ev��Y�A�Q�y��$�a�3��H���=�;ѷ ʩ�F��_M�_�#� �7"i
����ݛ��M���.���vŨ�&��kT'h��}ncv&9�vῴ¹�}�%���y�W�Ӯj����v�{(׵9L�K���`ͽ��zv�p�$Ĝ}�ₜ��Bo�L��x�KeS8v�ir����ǻ狶/7��xG_���� �Z����\�R���Ŷų�q�''���Z��k��=s��c�����]'[is9�^^�C��C��X��4YMt���u�l��nI�fuv�-��>Ǭ5f,;[g<<��.��7�_ݡ.��NN2yك�����=��q��J��B�j�yz�|HP�L�p=q�M˅\���$ͷ����Z�C���uY��l����q�g�d���ȴrWX��&�s�v+m��i��;�.��V�����]X��\٘7N0�%�a�ۣ��lFD�Bor�U�u�����k��ws�qX�ێav���n�ŉ���G�1!���s���g�����f7���n�.']�7��g!nӆ7aݪ�8���qX��p<�;��m�7,��\����l1�V��{>n�9��=�v3�r�pz�0��/olۮ�4����s��f]����:L`��w]|�Q��l��4ąVȋ ]���ҷ�wc��|�ɞ˹qr��w�==�/n�e�rg:8|�{z�7X�M�.�8�-��Ի<v䀢��燣@9��~����檱k�WI�`��p��a�T仹�g<��W����:x۔݉��|������a��:g7��؂z�^�7cY|�D�D��}���zk��+'sS�c��Fv�H�(��;Eh��i����{N��+K�����yYDPp�[b�"��n���+���ʶ]z��]����3t��O&��������n��U[
U�?`�3NCTa�w�]Ğ>>�?1��^�߰��f�P�83�j�HE��1�Ԍ�ƚ~<;.�'�\�4��蜡�n�ҼFo`U/w6FIO����3�z�����%�nT=����Ɔ��ْ�{�I�N���i)�Tm�v
R�@n��fs�Ɏ.���45%����jx�y��z.��; ��VZ�kEd����q�m�&b�T�Q�I��Y��\���dN��j`�ї�:0n������Z����H��O�����m�u�p4ۜltn1�a��TU�Kq]�|g�\��+y� �\�Z$남��ٶ�t�Of�Hs���d&8�N5Ӹ`�]���گ�	GPk�]3D�f�bx�Y]N#y�/�l4S�ćr>g�_�����ryt}Ɂ���PN#y�α�=o{^y�]GD�%�����ۛ�3�1{?E��,<�L� $@��1�@�{e�J7���8����"���������5���YQ�H�u�\N����Ƀ%4��y�t�<��X����fq�j{ʲE�s�i�$�Ļ���Ejd!v&ǯ[�a�9��t���<��W����m*�����z�Ԝ���>���U)���F���GƵu�!�%�%�_aFYuVqt}�5���̓�+�����>���ģRm2HF(چ��Q������[8��׭(?ʋb�97��nw/�!�q<����$��~��;H�D�(�o�������`#ގ�je �膦��p�JN�x��Mg��9| ����ołICǣ����ɵ�@]g�5^w����<��-x��D�*gE��H��Aw�3E�({��m�����q���Y�9�Zn�����S�Z�j��Iez����n.
��,'H��Y��WV-n��x�C��Ц�ӿ_��2^#�1��Ouݓw�H�&���˹7��a5���<GH@�y�]Wu�'��W�(/�j���1x��ʾ���W|���7y�1�4F��NI�o���&͚�"e_�*NP�3��z��M��N(�>1���$i@by��/[�:R��b����f�����gE�()ߗ���2j]1w���0F%�0����ܛ��9L���auu�0���U��M��ć�i{�H�8x�y;�1�[˹7�u��js��%��.mŹ�Zɠ�>̩ځ�0�b�U�4苬����j���ؗS˳�jZ-3L^��z�xų�ܙ���]ݩ.*N#Sְ��2��]\���D�0���==UD�ntY�!���V1i�]���1|�'I���q;�1�[˹7b���^�X���q
�����
��ìA��1`�9{�s�Y�9�XFR�ڛ����P�YN��ݡ/���Y�X~�����{�y�(�-y[6&�m��(@�U4[��)�s{RZc�Y��'�X�3��<����0�%����E~�
�����{�Nu����"��l-�R�OY����t@�{�4%���x$��ؗ�0jMHxth��3�co8���;��Bk1�r�P�`a��]�Ĩ�HĘ��{�߅3�U���N#�u��C�X5:�YC<󌻗v<�$������-Ռ�x��fa�Vs�Z�j�=ސ�t�	���[��s�����[���It��f�J�!�ω��<$�U%	���ʇ�ҩ���ՙL�X�ť�9Q{�x>����k�s؁.���:�F���3�8��ݸsz�`��s�6�tb�]��\�=m���(�OTu]��Rvw�z[���Z�ݻ&�^0�.G�:��޹����zvwlM/g��� �q���e"c�T�W��z� BrA��glJ!Gv��ZLb��#b���~��{F�θjw9�]���B�����fx�[Wskh ��x������Ø�d7��ǆ�z�bX��f�}�m��U�'�Y
��x��9�j�w�w!�x5:�1�홢�1{�j�3�J���>� rT`(���8g�De^0(��G��[�@/$G8DH�����f3=�"Y�ynb�� 24�|�����`�a�n}Dx���J�1�S�pa�LC�y�.�O��6u������u�>����XF�<IcҸ-++���ߪHy�Y�{�9��
�=y������;:��S�� _W�^���Lk��~fS��Q�I3?�?����mągw��� bf�;� U��4�0h"t�TK�c0+bm8H���_�p����<S,��u�s�z���K���um3�}��r�����H�9���q�E��\�1�Y��!�%ĆI�w�7��Β�������=�}Zh6w�o,k�6]`q/�)�q�������fS����ԧ"p�bnZ8���֘\=�����><�;JC�pfS��BSǘ;��� }ـ�R(�fD������y��JC}����g]\V=��m�^#'�ܣ�O��^� ��Ү���T���9x��B�V�va:иpмѪ�T��#j�#S�B�#9�!4	(Xa�K��]'�j��Ą�G́�T|��1c�S(��lKLZ(g���������$%E��ř�O��A\�~�hy�s�����d��y��0���C�ѐ�2�����d��lKD��g�|G��VKp���uv���#�)���Z�ͱ�����4Y�����gc���c��s��h�n7a�XL�F���qu8��t�b*�_@@~�y�U�E�xY<�Q�ҚӍsؐ�f�bR5��o�Y^(�w�o��V9t�.}�1t^�"2��E�.�j|&�u�Q5~�X0f�M��vU!�=�c�?v�����]�L�ȏl ��F`�!)U�2#i�D�f`��+~�X�C�z'�=\1�;�Yu��1�8�4��G�k#N��P�/q)�O�x�q*��ӊɅ�
(��
�:�D��H�zKe������{���)n���b�I��5�-5�{�z�c�VAp�/��->XA$�6[_[�3b�;j|8 |�z���?���|Hߋ����`��pU������� �{fh��b�����j��}��y�����<��"��z xP�%����2kYֱ��q>{߼m1NoA�lǨ�@��|��M����F�:}�*n�Н�����&���[�6s�BU,��n���{SXE�
''��F�U�Ʌ�$����u�zv%v�v�z��dӑ^�F��u��<rx���F`����}��6����u�Т���|#�\۪�۴ۮ����r[U҇�V�[6.N��W�?��b�[���E�y�I��nMQ��vp\�E�w�}I��l�U T'Z�ZX*�%���$%HcЬ�ѡd�c�ٚb��8������[�p\=��{�7,�c�w��v�ҏ8���HJI!�������y24 @O���x�rU�C��1QC9�w���f#38�������yz��O�xݯ��b�1#��z�����\v*d�a��]ךb��~�(��ꃛ���y4��%$�� �O���I���_K��!�}�2v�j�gK�Yێ�9īۺ�ն��=���1��C1�?o�� ��	��!�x�\&�j*d�~��������%*�q�d?�f@��4�r�n�I�f,����z�q��`�CӐ��p��3��^���E�!D��hI_Z�@��9bCƍ�g�K���ʲL��ɷg�,�b!�/|�]E[���ƫ��h�-2�ؖ���F$�,��{���r<���]%���V��Kf_~�m�慝v*dAN(����IS=��d�dt|O�C��I%� ��S4jG�����|�W�Ǚ����AlI$�%�;iUGx$[ml����W׼�5����WLbI�<����ݾ��ŷ�qG����>7�{ڏ=�t.�.F���\S_[P�f> ���Y�,�"N@W� 3�G��0y����[�d������w��MP�Zk%"�*��X���KJ��l�U���&�co�
G�6/&��D�gP$#7q�~���w�Uj�%��]V��I.���>�|��1��g���^���8Y��Z�gz;�Nj���˖�΅�lT��.^^���]2�Ŋ�a�%GH��k�w���Ӭmӝ=Rr�IDV���˻�1k*":D��sK�Z����#b����K,B�2�E��Vį��9��tR���'�����u�Cz+[1q:�mVqF���[���qI�~����a�a��=;Ԩ�Eֆ��	��9��.����2F�Y�#+�#ܬx��5�2`#��2�d;Rj;>�s�D];4yfq��unA2�q�f)�Ǜ]�������_Y�[�p'X��X4.`�y9�'#LO��㶗�w`�s1ݵ=\���UYl��~:���zo�z��ۡ=`P�l�c/b~BE������^1�Ǥ/��TMP�Ș���\׸K=�5\��tS��wS4��Iv�.G�K�/ �a��i7y<���$����y%\����m0�]��sL>������9�4�wqչ��ts^�C�����+(����~A�&����+ZR��P����o���H�u=N:;}�3:{9g�F��Fe�F�B������j˘�Q-��H:�'xm�̼�;6$�:�C��A$��֡nw!ܸ�{-��ġ��XV�82;Q��-+ت5����Δ��E�jW�3�Nep��y�;r ���{��zFm��mx����Jz�^��St=�O	�x٩�ٕ�f���'���&#��}��ޮ�E��P׋�X`2���*;#�N �'�8��J�Ah֟������{�e����/�e	u.�L�񉤗�b�x{��Mq+����ު��v=�U�����}������������"���Npų���K�q? �|�v� �H:7'f6��q��{��k|�4Vɀnxb�P��]����/:�S)���`��L�yz\�1��������Y��8�uߺ�e�]�V/7�r���o|���f���ļ�q�Pt$��>{���4�ṹ1��Pvʜ��Mǽ�{�����#ﾉ�R�~�1�Wmmb�G�X �������N�G&ب�i�
�i?�bMEi��6�Z�s�����
"���8.JD���bO��Ÿz��sE��!�>����(UdxX�:��h�ۛ�G��r!/"3�s�o�v-٢�ZQ�X�~��׌���E����>y3��>l���+�;���	s�����917��$�.�O���X�d@���f�4����k3��~������(K�s�J,Y���:j�bI�s�&d�J#���o3�O�dt���\1����d4ϳ��b��T<�9z�%w�I'��w⓵θ�x����i��!�v��v�`����3'O��{��̀4�yִ��X���c��*�Q;��c�ILK������� ���!���ҊhCV��T�����J���s�%<.��4��ܽT�\�s�pmOJ�ۍ��+vWq�V�
���y#����1���f2��H��ŭ%��� 8�V3�R	i���k��B����Gt�0��� `�b���i��$ZW���E�_�K4����bԖf�>��C4Y�~�O��=WKmWZK÷�ǋ	J��|hJR�Q��ūwb�խX8=�u��h���x����b�?6����G�a��Rx�ff)�,@��>���+r�~1t�?L�d��P���s������oI�1.
G�ē�����
�n)j��Lq�
�Db/�����ɝ�d�q�I�1�1�X�{��8H1t��(=�����l	�~�����!��8������]_�P*�����ѽ��>�pE��:tY'B�B���&eB�O�po f:ƍ�wlݦ�Í4)�D�pS�IbP^P��q����̦%�>�uG�v4uϞ��}�a�A�q���sO#S��&�7�)�b�b���k�bof]�}�|�uEe.�n{�9�"�Q��8��1��d�:=6}��4^��x��x�b��Y����Rl��ߟ:��3g��q�=�{Ч-<C�u�컇r�~�����캱��C:%O�i��f#_u�eI�m�|z���f�(�xz�4�5�z���<^�����������3(2$�����[ot�	���ɇ���7�� �J�/�K�~Q�يF�I��"���v% ���!� gLR����yf����$�c��RZ'������k*���"fX�Ym���k}���q(�ϻ1i��^�g�)FB�6��~ԔX�x�x����V��y�޸�S�d!�nz3���N�W�﻾��<O��2����A)M,[�S��ۨ�_x	�Q���enG�8�&�0�:Y��:q(�P��Vs�qǹ���:��<ICd�xx��~H/��F[�N��)���ڨ� ��dxx��n/&fb7�8O��F��� ���}�D�F/���+��DP��P������w~7��+������lϑ���D���C�?#��T&}~́N!nQ��u�@� ��=S�q���W�j(����Ix�ג�y��C�W��<<�&�S�K��1ud�|�&|)d�F�Q��ЊPV)T��qQ$�t�-��䦱8�w؇�����S����.7G�b(�1 �0l�������mo�G��K����x��c����~���wֳ4��O�����D9�g��#�����L�`��L�sƞ$�;R��u�5����N�ތsYƴ���e�U��=\�'yۧ��{�y�}���E�j��m�f����}WUֹ�R��#�8
������� �̃�
� hx�[9�C���=^�0���nh�;+�n�\&���\睹n���^��F�y��F'F5��h�qs ����ӷ�:��s�]�<��70?\w��S�c�Vv�&��D��2��c�t��4Ů94�#���ʙ��q;��\DJPV4+X�VD@�%��8��x�۹3{�x����{�ǝu�/�f�Y�x4�{�{ƽJG�����G�pj;�~{���=����9ޝ�i!,������^C�A~����4�j!�C��٘KobeR��2	-ç_x|< zfU�L����S���1��^y-�R���k̯2x�Y�%Ty�y�(��F�}�u�y���D<gR��塚�)t�3.��B${kkےM�̨WU�'IU+�q�;�������=��m�	f�2q�Ҟ]�z���I�����̑�g*(�^�����f2�BCk�����x���f;8s�zQ��!ju��$�Hc�D&��y��#��6Ú� � ~�R��-�T3^T�w��!�Ǖ��uUԠ�������^3��I��!�?�|���G�FGw��"O��FrApP��EOޏ{�:�HDf����(����>� �S	w�YI���g9��u��qQ��P�^��ޣsԙ�j�LP[�S4��K���_������G��ͻ7;���w˞���//}>Kgn߿$�%��d��>��E� ���O��(�.�E�t�<0j�Iz�oq���w��1��=���������Q�|����-2N��I�1�w����LOӊZjЁY0,�7/����Q3E�s������<D�ӢV���q��n�����e݁���l��*��I ����bm����k�QI�
o�,�����jh ��-l^.����n�t�v�w7��x=2%�d�����s��՞�����X��l"�1IDJ�qDA�aW�,Q�`h`QX�Q
�Ɉ�/�����1���t���*\�0�xO����R�[j�����f>j1�4�5I}��V�z���^k�tUl�Ɲ�N
����2�H�u1�;33q�y{�蓱T~�"]�2�Z��a���2S�!��ج�z�7��^y$�ƶ���by%���Fъ��C�rF�O�bz����y}�R48r��2!�\�WW��oww���ů"��B�A�v�E����Lj�4E8�t���U0��K�t�������w�O}ऀ�J��+&`C���o�#�+H�&7><���������Y�;��{�Rõ/� ���>Y�A����G���u'��>�U\�ߵ �(J[�L� &<9�Q-��88��(.9�v&dfB,�{_��t89���b�֞�O<���֒�>�v!�n5��~��`�>x�O׵��������ī�J&�6s/��6���-����o��dΩ3W�lg�ǋ��h���3ƴFOe����"�L�,{�����{�dE�Oh�8�-U�Ύ�X �S}�f���F���5�Q��kO��w���f�u�����W��q�����զ��:��te]�r�Y�ޔ1�8�^�:)���/241f���kw;ۯhv�qmU�]QiT�9�����;f�\~&��?G��߶aF�vu5��οsٷVr���o�{�B�������r|χ��oC�ʕӹ<�=&7�"M7��N����6Mhɳ�Jm����u�������[���F`�NC���j��+\��g;�5H�4,^^��k�S��E���r`8ӝ��z�y��7�wD�j�&.n�n
r�;K��;{Sb��z����V�<�G-`9z��-v�w�e�]��`��H����*��y��,��sn���֕��V^�)vu�l�μ:���k�vv�^����q�nG8�k�v�up��nP�j�y��q�G��f�f��K��ދ��\�\;���]��{���݇�<M�>�tݹ6��ɭ=�/g�=��wk��k��M��E��=����Z�ݬ����u�q�Gx;/X�D��b��e�t=�w<n���#��Q���G���L������14m��������W�/Pnx����[�u㍝V�gB���R��-��u>2��*�(�&ӦECP�2�99��]gθ;y7k3�Y�4$�=�k!s�TpiN'
c7O����n�9����9��z�l�9���Y�s��G��6'�[
v<ع�U���,t]vF�VC���Gl�d'�u�i}�
�M����k��nzkZ�N�Ç. q\u� �ݟ�3	���R���7�t�"���9��]��A��C�X����(�5�0�+:f>q�
ly^k#ټ�F�/yѝ��W��$����]x�8���#��3b�xvM78�I�5|O���OL�.��y���Ѽ.<��mzqhJ��ȝ-��.kN�4��N۫<kgה��<��ͭ�v{�����T�{F���5��znqv=|����yu!��`C�^����t�^����n݊���F��g�K��]弉��U���X5���v�<eh��'�Px��v���5[.�o%ܓWL��� Y_rY�'���$�_����#�mO�k�@�d+���`���e#drxOH�Wi���hy�U��\d���l�����o�̏'����t�E��C�[���Y�}�|��Wq��u�;���ÓF6'J`�IrX��ͽo+���s��B���K��<)�R������
k:9�p!�����۩�X2Z�Q+��͗�pm��du��l�����v��vu��riQ����M��{��؎�*��[�H��4oJ�ɱ��T6_X��ʙw.���o�^,����M���#,N�B,[#5F�9�<�����Z��w2,A{��jؼS�Z�����{�(@�i@���1�kγ�;�����:O��3�v>D'wi�sw|X,_v�y!����8�������8�U�{�4swD�-�8m	=qs=Y8]�O�|Sŉ����{A�d�a���l�^T�wJ#K����UH++���󼓽��r4�>��Z(���<&[H}�ו�Izu)IP�y�e!9�s���*l��\���j�^�{D6��-o=��A$2�yCd�[���0�ftZf�RH�m��a��41��VM��ie�}�s��w�	����ݏ[����q�����Mx.�n��$߼�������@�!Q��6�,�� Nj���g�UDf)�� s�޹Z�ց�m��)2�n�)lB���Į��*h���{m�	ڬ�G�0j,�@*��]��=��}-�X�G�=�������S��]�|���q2t�T�`�/S�? W��${:������P��UC�}]\|'k�V-��6T&IP��dȟE��U[F���@?,J���g;�=�w��zB���پ�\�1#����q��&g}���d�[��>ؗ
�#j!o��x�zs�M�V��z��~As�d-Y
�&�r���"tf:�ر�=(��e���I��G��<M#� �����PْoP�p���.��=�">>����FI �,���Q7���D�Q� w���7� ?�o,u�K��]�;񭏫Ư�o">�6�g�(�ᘿ��ɟ�c�1�;�<O��V�����x�+
�X�~�ڍ�8��f,���p�YP!)[z��;��M,�ђ�xT�{�뢲��܄zӉt�nI`��{ŊVև҅9�֣����!b�_��>��{S���4��_x }�	'mD��L�+<��{K0An)
X�i�\������6�cM���p�縐�(%���s[�#,s��1-�j��c��J�w�;�>��[�]7��}�3�/��V��)o�ԍ��1�!=7��0M�~�Y�62�ux$/�	��DycjI$��qAnȚ�]�]�v�SyJ�x��e�^{Z���˃�X|N�]GF��p���u+��/m<�z�.�k��AS�xs�a3p�ʺ��bR�8�x�L�7N�ۍ����ƀ��Q�9e ��ki�	��|﯄F��wPc�sr�J�h�ƅ- ��,�G���5�Aj�l�� �{�QK�h+P!�p?y�*�)�{������fi���)"?�ٿ~��\�z��%=��\�~�`�_�����RF,���?x����Nk��<��}�;��𹳸��R=1�Øz��s�Z5Ha@x�,�&%�2/>1E}�� �l�g����M}���-����mZ�5�����������o�;,*�$��.2�'PN�T�cJ�(��0t��MpOPA�@U�pǂ��mM�nI����^��~'����e7�s��D����)X��lD6����(xX������!$���k=]�6A1�����}�w�*WF�2�{��1[�\7h�@�3��rN�SvGm���f=��Q�����w�{·dFY#E|��I凼;ޘ�4�b�N,��o_�H��t->�{����EP��ut�>r���=��\���7׽f�:F�8ARe�6UT�۴�E��R�i�bl����A$��H�4SQ��ܙ�i�^��5����8�Ƥ{�	 ����v�
<(�5��s+����LJ��MsN��;�� �e��5
D6��VYb-���Er2U�Y�#Q��������X�G������_g�D*@�È2o����9�'5`�xxLW�;�hcz�{'9�}Ľœ��7��8�G����͐o�[��Cg�;��5�cv�]{\�km�iE�U��k�}��b�[�5UP���6�3��07�f�#�#D*�T�Ҋ* _�v����N���i�x��|�Ka��=��4>�nQ�dVR�hة0w@C�H�VX�����M2��8~AR_}�O> R���$i��M���]L����� '�~@����?}b8�{��ų���w��#�$�}Š �{�;�G ���$p�]�p�����I�����ƾ_e7�&�[���v9��n��0��1���+�	������[�}�YgN�*I"G��6�C��ku틱��x�妐g[��Xm��J�[�Aeϱ��\6ۜe�G9�x�����rC��b��ݷ��v�s�m&�	�q���u���ty�w3�b�hx�&-@H��"�l��Aȶ�<��r�giz��2t���}W���3�n� ���m�$VJ��e,ŭ]��������=��~6-(~� g����+y��v���S���O��Y=��3��M�l�6l|�m�lOp��+K/���,��7��MYã�G���J���?}��/=�=��	]��Q���ݐj�8��B|�I˱51����_oM_V<Kjl��y��2D��7xyߢ����;��ѓ�~���&K0+,�<��,�ry�$z�Hn/y�z�ւԂD`i趼Z1F��`�m1R�O)��*cɲK��z��ĎG�]�I�}�ub�~�_�8	���<!�X�S�Y�+��Il��u}���ڳ_��XbŢ��$N�&57޿1!bW\�����3K�nN����#��І9 !�B4K\U��X�ZTZ�te����$v�,��}5��R�Bi��q&�����	��y�<ILo��10�)b֝�A�q�;�#�iY�� �+��6������¬=��PAxb���x�n2����u���}��tQ��ww��n�1�Cv���0b���ܩ���W��K�8����Ƨ��iT��<��e�Z��vyД�^U�	�ΖtD�&'U�[W5F�|�*O�)��m�,�q=��.�6�"��'���ܚg:�����ee.�4M�;�.��|t�"�'<|�o~���9��v�����u®�^,K<�Ԡ�������������>I�3�k�)!a4�5IJ����l\\�,ͰI�1H��Sӳq��$�n6�S��*��-�b�n����m��lDV��B�qs)I��.ln�j^1<V�O*�������]���ҭ޲jt����U���Z��\��=r;�'�c76r�	un���WP��1:s9N�U�ܺ�4b̷����w���ɫ8MV�!<�H���)�1L��6Du� !����x�&W�Ӝ̞*���t�#�`�]���Ҏ��&^_k�'z��v]�/�(8��W7	G�PǓ��l�0=ŜތW��O=�{�,mla�LJv��̻9�z�9�:)���_�jp3e�+��N������=ss���{N^G��$1�]彗����}tw�]Wy��ex_������-��l��<���a�V˸6�킾,@1w���b xٻ�tI��=3��O��mk�;��!�=��>�����#=5�M^�Í!�r�v���7X=�o��0��="w�����?��0��kX;A�������
�2e�ܻ1{E`�hz�J����v8]]�M_C����2�*A*���5S��sZ$#����Y=�x��)��k*�
y��پ�O3{���	�o3X�V���̷M.0{Ç��ٗ��[�	����~��ӕ��*���e��Z�
`���Q2�3ҫUM[X�����O�Ĵ�����/kqJ�c�� D	+56���Q���/���@��DU�h{�v��_X5d�pN����|EFxX�=Q�&�9�wl5��%
��:6��������q��.�̂�rp[�R�@TS֩c�]�px
@U:h�%���^?W����c|��˙?|���x�GG?O�n�v:Mg���M��b�+��}AvC里/q-�}"�<�������z�����'��,J���~K̸uK���SZ��z��@��ծƶ� =���kUI'�`�ݪk>ޒ�E�}
�+1��x<��}�̓+�m��=�z�Cv�Ln���!vt	�ٽ�%F\���Y���+�Żz�k�vo�u1ց������q�sx�^��,�x����N�UMU��A�bt�BEULl�<i����A%�MN�ַZo[F��=�U��v������G��dR�X���������ڌ�ֺ'Zb�W|&�� �j6��Mm
Se������:٬�{��ݜ��N{�k�IHj�+Ҏ���� �|jo��4xT³�}�he�i����2~ "���	)��f�xS{�i�MF/u��v�՚��oZ�����������w�~M������ y��Q1�o�(���K�B�{�^ea�]��QG�����\�T!KfET"� R�*hh�RA����e�x����SMup��2���h�Ȃ�N5K���N�?|��
!�U1]��.�P��mvϭ��Z
�lsoP[��x���m�T�bTj�Ph�ח^��+`�?d�1�QZ���bԶq���!�0g� �Z<7�>��%$�b$٣h��!���BŁ�X7`��+�ǧ�_z=��QEtImW�>+�!t"��5��$d	H�:H�l8����H.7mf�Ѻp���c��RK�w���i���A�E����߼j�������Ʃ��q��e�lu_شdM��W.��9pU,�����;���+���{l��;�����/�5KrZ���m�J��{��d� ������?)`z:��DB&����3��8�=�Dwiy�;'�D��J\���]k���ݾW�Hn`;b�~�]���~�µ@�������3f_͍������a��#����֙"/��p�N{�Fo�Ť~* Y����ؽ��нUQ�����U)���0��>��m�I�{=�=4��5�����RT�ᨋ� \?.o;�N�?g�sb�}�>�FZ�m������}(�Pk��<���Q��kJ^x&��֥����f��-jw���������B��s�CԞ�-��e>��qb�C�$} �&Whm�p�,�D���qs�V59{�����1�H�(
av1��¶d�B�<>���c/E�W�k��'H��±����#)sɚ�)�H�"������Ѡ��ʗn�6�/][4Y����qx8x���^�m�Ƌujv'n��k�e�l=�vy�8܇=E�^F�7:�n{nq�)��[��\�JZcq��li�W��s�QCn�-5�7+�";��i$E�*��I�������~ֵ�	)q��Ɩn�4��^�ځ/�DɕЦ�ߗ���z���'��{���.�w��S4�50"��84�������铻Y��N}H��A�bN}p{�-����9�b�!(|�0�H7r���BNAu�k���n/�0�6~؀O�x{�1�͜ϸB���$]�_ą���ź/m�
D�UU
�f_���^E��T��x��x�lrE��P�<ڮu�0��ग�[P�3e�Ss? R�%�|B�!��獵O6��}7��B,�q�a�2���P��(ʘޙ��_M�kzս�� ���|�؛8�g-��A�y�o�bn�P���;+�����3���n��o[/�Je��/�{�g6M��a��!1ɽ G�](;�6�Sy�K.��X�)�M&$����G]ξ�Y~�b�D�e��
.���*rҁ{��8����3���nJ�cDx m�'�%AD��R,����Vh�FU�2T�aB�<�V�A��'w<`h��tD)���VL��>/���{�D��8�0&�ad��v�<��t�����������|���d� n��!��_l>����m}M����
�T��2���f*b��m*1�Ϋ�dv�d�� Z��=�>N2�A���~�U��\��Rc�}"�T��gs[]�*�:���o2G��F��ڼ��L��#>i�;�U)�8��A��B��5� %��N�:fR���e��;+�,ߩ�N|����l��3)��D�pR���)d�(�����^D=�7}.�<�?)��}�!��{ȣ׷��wߓ�r(�wc��\1�l��zk�"y��@5o5�������_�ߙ`ê_F�� �į�s[N��s��	��yWS���7�m�3mڳ�v+��Xy:ˆ����3��@)��(M$ٝ&�i�e��#ܥ��l*{���݃ǳ��;_��cZ�j�܈��o)W��x�A�Ϧ�ړ��A�I�rK�ބ"��@��L������"#Wv�
�[�<,����ѕ��veٮ�hD�
ɖ�.Y����{��e�NqWb�9��[����g:��l�(���a�R���.�]�7�gx�ؘ8�O���zH�.���ݷ�H��˗�Tb���h�F��LuwT���9�I"8��	�M��E�<�����g▽|�tw����]s�e�Xv��臖�=��u�dZ�����c�X�P���������:¢�7���е=Y٣Ktt�ۋg�2g���h�\Fa�l~���J�v�#%���:w�DO��~��q�=9�U����yƬ�us6���|�۝�^U�\��e���uj��>�ͭ�gX�� ܰ�m��`l�u�{���q�q��rn�k�:6�u�iˣ6�-��B�u�����e�����òu�g�X�z�d7&�!C�s���e��Ũ͞$%��DQ\�m�[2�f5���]9��H7L�m�׊�gwaݮ:���[���h8�g+P�q�
7���wA:a��t�:�U�(�j��#"�ba�.�N�uʖ��m�ظ�%��h���v9�.띳gq�1)�4�қoV� x+��'>�9n�[��2ŭ�9�js*�v�Gas7�۱=	�5��h��mD��d^�g�t�_����^C�P�����޼([j�,Ƕ��GV�����UR�e�a.��+ۯO,�l����Nyv��re^.�H�{�����<EsX��7�:���uc/S��k�XL�pq�;�
�q��voR�d6���v������j�U���x֌ܙ�zۗ�,��\��c7^Mrܜvtx�t����0t��%/EҬ� ��|cN�έ�bML\)Oc*��A�=���a"ڊY=�	IkK��4�g��8y{���vɚ�� �//	��͈��,�^��,��f+��,�\TT���dV�z��B�!"���b���"����v�/wS�9����|w�L���Vu�'�2Z�=��c��{ޕ��uh;\�z�_���^�m$0��s��3�wh��@����(̐��xP�mZ&�������Oj`7�%��r��D��tt(M�x���Y��Z�7���x)�����4���]ٳ˟Ι����8���-��X=�?����4K��H��K���:�´#�}4�y�����_�zh;��gLQ�潚=C��{V����(��zs��v.����7�L񞓨K�X��pE�:�Ů��5�j��ǉj���P��E��f�pm�g;j��]����,v�ۦ,�e��]�`-��Q݋s0.탨8� rcu��v0����5ٖ�Wsr*\қ����{�d��87��8'��lcq��\C�8��<�jL�u���˻�����������z�]Y���Y��3�"$(�N��<=�s�fc�11�����6���CADBp�@�����5�k��3MD��ʘ���ZE8-�f��������pj�3�ܾ�3�H�]	0�H�ؗy˧�o|�fjh���m�p�T6�����烍�N�[�}���O^����T��bK���jUDh��ü)b�wN��j�V�фWFϞyً� I����	����Φ)�}(i��6��L�@�zR.Դ�.i�&7�EQ3�%šw����_3�ɭ�z�v��x��8s��b,������@�t)H�]���n.>]3E�9_6~U�{�g���(%r:���9:t����N��{;~����}��jL|=T&��4�w����f �-�� Lj�O2 ��1�a�IH���I}�'s��U'� �t�7���FMT-A(��p���i�!'1c$מ�(�5�U�h�mZ��C:�cJ� K���Q ���I	�����y�w���=YW�f�붻9�ܶ٥�����_]�UIY�X ���Zl53t����e��hݹ 
6X����ɴ�[i}�	��fc�5ŷ�u�}U���-�m�e�U�3��O�r<J�..#�M8�Fg@�e�;}U5�3�4�,����A�ߢn��&T���yީ�R#�O9��3�H�k�_�zzv�%f��3A�@�-1��m���&J���LL ��S�(�EM�)�*ѱ8#}�
��W�Ј_{ϥ��	�����ud��vo���ڼX���c]��+P1Tz�y��9�͸�\�r��ē����b��C�����(�o;�1Y;�&��yYY��*����#��kn���ߵ���Č�l�O�X�T��'>tDg�ψ��"M$o�ҩQ
Q��s����W]L��Zf�b�]k	�=U,kU9��3�2(�b����������ʖ{bp�`6|n֯m��:دn��B�:��ksp]�i��W	���2Y���^$��m�#�K�nN	��y4��6^�ǌ5�^�Xv3��R��v^���2���N\������(�»h���=�m��d���3(�E��3�8�|[����G8mbM�+t1�"�R� ���57;<!4�O�cZ�s�i�����N���? *"�B?B��(yy���j��m���T^K9jI>�m#;�]�(�T��U���%G�iu�[�)���������b��O�h��h����1�v�(ڣ#���j�x�=v�p	��;��	��m���e�*'��tFġ����i_֝��l�*L=}���;!s��"ϲ�߲"�r���êD�����c�#F
3J�n���^|N6�O�,k�|��e&�8�ߓ�/�}�*������9A��lExq��9�B�	D5c�|��қ�үFub�q����IeM���/gk�,(�(����<�ï���-��\���I*��=}��4�)x |͎֐XYfs">��������у��_���*�0 _B���jn8��$��&*���c}����d�$�2D/���v��ё	0@������R�B�o�((��{[ia�Z�j�]n3�b�KAfN�F��X���H�>��?aul�\r��㛕�\�܅va�+Z�D���֜o��A�}�cL���|")#�Z; �>5���"����i#��.Rc
'���@� %�Vc�ݍ��r62ѫF��Te�9�G��f}3���	���A޷�Sɚ@�HIA���\�ѪH4��Ш�y"N(�D6��Q��Q/A)��T�cg�yi�s��_XN,����@m�ց�n�B[�$tg+�7����y�R��.fQ:<56��fV|�����	D(S�e��_L��Qy�L����/�-զڑ�mv}3Ϋ���G�^�(�zߋow��x����ּY�[Q��aEA�����-�s��E�ыy>�w�C�{~pD)��E�U<#B�׋}�T�M���$�qB(�����Gs;�F�u�ˤ��ڳ���4 	cɺ�Җ|$v����7�]�;+\n9�����s�Gm�����7�'Cݝ��*\��X3ֽ=��р���I�H�-{+�����CO�E4[@ӂ��U�YIy,ݰt����gg�M�\�f���Ϳbվ;ߟ|v��Zw�kr �E� J��K!& On7i`�MY�C�R�U��.���>,�M�zd���=��G�KN=j?��v�%��}���Y AMb:͒��Ԁ:�U�ۂ��Z����t�����]���R&�$�{�Ȗ�ξU�;�����D�Ʌ�yF�3n��Һy͌64�G�W!F���Fɐ巄��뵶}����z)k���G�x�;��������'��˹:I��u�p������QFֵ�b<��{y��8|UJ�%��QP�s<Jp�m>��/r���,�_{��W�ݍ�C�v�զ�Dۍ�j�A5�k��;d#��n��5�����1�U)/���t�7�w�D����9=��W��c3^��ꋦ��Z�g���'������;�q����əfn�
OC�u�iK;Ǻ*�篶�Z˞P���p�f]�"�������5�+2.�A��ٸ�w_3�����1�;�$j�9��r�i���a�o�1�BL��' YnF^^�	r��{����s��9Z�&o�C����$D!�u�����J66pH��&�ж.º��{�c4,�{ٰv1-������z��0v퉌Q�]���^��#b��Ǐd����3Z��?{R��&��ۃ�������o �����k"�5)������ݟ���Kؚ�Y��3/0�_r�"z��'6���H��fc+!@��>���==QuP�&��K켋�����"1m�(���L-�ME���������{�ßŸ"�ޠ���������N���P5�vy��''��*)3˻�_�����{�<(�svv絴�P�ͫ>�b����4R��W3���.S��-ﻗu��Ѱ���M��kDɡ�<�j�r�ӭb]\9��*v�s��1[����f�ѫ�{�}<�=���o�]�1�������ztV��v��0�F��S� ��ٸ�K�7��
�����/��Y�B�"�/��|3�-];�.�t�^h&ͧ�¿Eܺt>c\B���*z�}Eֱen3!ک��V�D+-k6��Qq.�u����t���N�չ�g��ӈ��m��F8ni_,�
S}+8�/��-��.�����$g�8����0�9N��ձ��6�Bu���˧%=�{m�d���Fр ��6B١T��xkE�d\Ъ5P����e�n���.��c�4��
!aF��U]�*7�2b�(��p:�m�q�(���T��bD1	U��iA�Ը+�:
�%�"�N��Zg� m�{��o�QA&�n�]��Xty��	Q�V�ʨ��"�����cd�(Ŵ��u��'��9���osi�LG<P}()��>ޗ;ąJ��j 	")�˹�I ��ϞZ�٢�zkt�����2+) ��G�=sMNG$��o�����?��t��6��D��J(����ٺἣ����6���N�w�ՙ920%��3&���zU�@�.TP	e�0�*"Nlqbn#|��3*�hw��˭��s�4����~�zX�X>D�шJmhe�Y��C~4�~�M��4�p;��)�P�wT������ѫqb� ,Q�t1-'��]R�}m�"0�M�� ��sƬ����!��ɋ���.	ܨ�NL.� �l���0�ʱ��5��:6�Pns�㗐��fm˂��r=�����;��a�c'��v��J�����gk���&�Ȇ�ja9)]i��s�V������8���n��쌶0�0� �Y���~���&E!�B�\K�	��1��G�ݱUqF���ڱ�x�m���r�9X��(�F"$0����w�ɻ�3��;������9
�� �������3L�b��yp0�+)\�9jM�YX���Y@j�c���w�~�\i��FҢ+�v"��vimM_�$mdoYcb�S���Ǧ�VD��:bf�rm�Li��`.$��<я'��	H�؎ȗ~s]�ȏi[c�	��ǧo;ޛ6rQBI^)��`Ζ*�٫(%[qU�Kv �f̊Ag���|ALaI�p�6�sO���iU��ov�����lq���N)D����M�+�*�z�̇���aa�Je6���{�TZ��vD^z!@�ܴ���zb�CW�Ҥ*1�Ƌ�	d!	U.�r$��\:J�qչC2���_UU���vf��jƯxDH�������^j��f3X�A c"x�lJ����g�A7G �bh��� �_2�&U�������}�󆪆j�z����[��_s������8R��]����W]%�'hL�ld#��g;ٟ}��}|��4lP�������7fA���;����  Q�=ݳ/{�DV)hݸk*�||Cn�aU���8ԅ��.��eu�U��rЩ��)Lt��CZ��8v^��*cU������p��>��U��= SR��ɍ9'�l�{\`����!��߳:�Y�~�u��W�â��Fܵ��3ٮ���s���A9�D]�D��̎��2c-�kbEa0�V�� PVQ���������"9�.*���u���81d�{�3fJQ��+7[���O����Ӭ��|Zm�9�l����P������!��W�iOFj�86@���r���7ٜ4EZ��P
R#
��oFnH���<��YDK�F��;<*��k�����s����j�m˙ɭ#�R���yF���z��]��.]��e�S�Ꝼ\���B���ў�����c;�\l*�7>����ݮ3[�3>ك8E�r.&�C]��͛�M֤�Ȝ�UFQ�&��\n-=�\Z2��=�ڸ.`�Kq:9�5Q��{�7^̒0h�H.pؚ��y�܎���=���}�N{u��o�U�

�W	�<n@�S=� ��쟌�>����sl��n*��!�K�|���v
H��6�J�(2�F�o��7��I�_z��0�w�O�w0��ͅK��ˋ�w��N(�Rm��������ۗ4�H��R�4o: &�������>�*��pτ�']�l�튣a�S���&�nN��<s���B�=�k37��ZNȀ�KD7X��1��1��?���c��sH!Ç?w���|��ʽ�,kxv�+#lej+1��paze��w�v>:�t"!�k��fV,i����>� ���G`BUI}|4D���|�f[�~�q�pEqQ���� ��G
ٝb3�V:������]�q��i��9� ;�&=g!�zbH>EJ��	İ�F)T�"!*�x-�Ò��}����8w�㷼������ћ"(�F���*� �����V~苵mo�W�?T5"���<�v��t�pl��9+�Zs����z��M}�쇈d����bc���bʘ[���ˌ�PF��5c��� �[�{�u}(�;��"��
=�h;'�R�#eJ��^�ގA�cg�X`fL���]�];&]๡v�&��=ț���i��f}ִ}����.�(�T��!&2�ЛJ��<<>�|^��ݟ�x����
�e$@���)+vRV�J1���t�-���~{UZ���gu~��������Υ�1dulM+�m|�j�K����L�V����� ���� ; U�i�u�a=dǉ��G ;h�}HwЈ�3X�jF�q4������w���be�e�����W�']��t�6�U��y����ͭ�{6]�gi`y�eQ����t�9>�n�ٛ/h�N��J܉}�P�SѮ�{,P��ER��/;6�r+1Dő��șᔅK
���Fm�w:�p۞���۬P�j��٥sȋ�!�X�Pkds�Y��~b�v�s��wu�x���O}��L���t��g4$+�SR�Egc�f+�vn�Ow�]�}�8L��;��7�ʲ�ν�}@ڐD���ꤒN3bj��l��&�s������v_	"i�b��%:�ʅ""q	5��U˺n��h��3KFe'���z�E��U5w��E�)�QxTE�m�s��]y�N>��*��2kk^%I;÷qt�&b|oosTv���ƺm^'֠��y�˨��:Χ`�
8�d"c]�[R&�fm�j�S�R�")�#��[)�P|^x��r�@=tv�ũ#n���nx�c����ӷ16�+��P����)�흶{�뛎c�Bu����i��8�s渞���{]1��n?t��t|��.�>z
�G�x�U�)�ce�����6.A뺜q.:O;�I�vz|On�!�:ڴڹ۠���sC�E���Y�\���9'Z���Yq���g=�Y�v�t:9�W0tXy�#�������m��uǕ�,-�5��a�C���sr�y����s�̀Si�]�'2��4���:�2u�g�M+ѣ��@�nS�L��29^�s���
�{��i��5�<�w*I�	��N���)�:�b.�oh�[sL��]Yg�v��ݻ:���ƻt��g�����¹�������F��^�̏K���*�Z�4��=qہ�v�$Hݺ��'�^�A��C�{�
��z�q�<u�׮�^ꚷ\��]v7�]�p�mv�۵����j�4s��9<��ڲ<�]4�'n6�)u�<s���x8�ݽ��\�v$����<ѶU��km��㶢\c���Y�N
�b����ϒg�c�2���O��O.a��K�<��Ց���s�b^ŐcI���~�W��fl��L�y ه�ھ��3W���k7�mZZ~���D	/&\�іPu��]�V_j��x�	w��?6������!����eH!�ۏ���������X�ϸӹ�=t�Y����s�J����U\��Nx�ae��^����ݘ�/4(h=}�+]��/G���<���y��r/r������=Y��ۄn)�/��(�l�1��n��K1;���O�|0����[���C��vspSqp��dy��{q��q�]�F�c��A�t^)\~�}֚Џ: ����&G|�{�������"Yü������ZN��$ap����&_;逷w�[������g^��}���b-v��a�p;�nU�R�9���uٺQ�#gHW1;��x's�;X2�:y�۪G������Ϙ�'���%�V��$�<pY��v˗pU��e�"�JO�Q���ۚ�^��qُwz^,R��o
E��&�����PTM�*B�1��"T�S팔B��i�t����3!_,�_�S�
Vy~g��Z<����R��V"M�݄L]�g8��_�ߠI����l�D ��8z=����� ��"���O�j��i�O�Z��Cy��KG�C����5\#�F�G!���+
o���۔e��������YJ#���؞�O]2r����x��z���**Md�>�t��v�S���z��n��t���Nr��0Ԡ�"�lb\��6��=I�_�I�v��hPaj#��~㽑>��"~��_^x5(eL6 l�ݷ~�3�6��Z�Ƴc���Cƕ�n�j|]pk�~�3s~i�Q�"؄m	9���44�.,�����=��f��}j5�6��ؘ��Ѣ��P]����`3<�NOC��˄k*�d�|����fe�.��(��\n)�RS⏺"]��hCT�S �:C;)��k Bi('��Y�#U{�Nd^� ��U��Ue���x^	s$�a���ۇX�<�mu�G8��,@�"�a��]���6��pۑ{�GJ�,z&�a���䛉�"�/���Sy0`":�/���u[�d�,��q0�A�,T��.���ڍ���.�5u���L0�r$�wH�����y�)� ��x�Ǎ�=&�4MF��s��j����|V*RQ�w�Z�y�F���N/�W�lpvZH	�2
¦*XZ(�HY@��o�=�KlLMWY�e�7Se����)̶�o'&什����Gɵ
I���'v��&��$a9 � BSc��9:9�,�(�Sy�I���\�`eQ���x9e�����^b�suΧ�q¡Xԫ���v0i�[X'�
qk�i�U6p������q��cy��Omκ�Aqa5�m׮ܷ&�9�d�]d�n۶wd�mvڐ�;�9������؁F�\{qGgE���r�0ۗS�ro=p�{TWfw(0����ʌ�s�ߟ��ۡ��V�B�P��R&�uA�rO#�D�u�Π\�l��B)A�go:ۧ��x��k�<i�k�����4tV�,d&�����9��f�OF���n��A���g<�f�#�nFj'G�o[5�	u���-�"MqȂ�$%��hqdUo9=y �B�߫%�ǉ�Y?�]We�Ae@d�@�JU�N/>�^y�>Y�����;�G�6D�i
�P��vo���f���%y5T+� ��~yf�Z|
p�Ӎ�^.܇ji��݉�l����=�Q���7GP�!d�n�w�����ݐC��u1~z,��ޫ�ϟ�o}쾻ޡ~Q3�#"@��=�-o)�͚���(X+@I@p�&ms��gi����Zk�f/{����V�����ڂ������B��޷��3f�F��p"N�k1�AlWGP�)��ie(z+E�N�M����>�Z���T�;�?q܁��BcQ�a��U��fr45vx�*��(�
W�����56�O�����2k	K�S��2ia�����PK�<$A5�%�D"�k<��Q��>�e6�	�hB���[;����)Z���;�
Bn&����*�Aﵿ�x����m�ﾎ"w!���́6(A��3�otY�=PI�l�0��c�p���|dr�3�ݻ�~"%��b����v�L�;X⡭n��b�Ч%��Ul����]ԙ5�2;̴f�f��.�������%�{$�J��������]s�kV^��O$E؀f�ٓx=-ɧr�o �.D�Rw��ʱb���w������|��kj?��f�lD&�����KT-����!�e:5�������}�.n� �ϣ�79�[�U�}yCW�����
��.�6�v�`�q֤\����}'٨j��{�\���߾�ـ�j
����FG/*ݓ6���"�F祫8���z�-9�h�;�z.s+g���̼��q>{�~��kaU��ֻ�4z�W�z�r���ȉlػm�I� �=Z/vG�7~y�����J��M�GJ�:��q�=e}N3͢�U��"��h�2Q�ЩS9dc�w�>�"�.~������l6fp,�G ���[�8k}�q���%��E,]�ī�����k�Z�EX<�P"�i��Z���T�[|< Tf�Oi�f#�څT����.����Bw3��}n��!R�h{Q�yr��n�=��x)L�P����[�B�]���_m
�{�Ti\a��l�k�v�9�
�X5W*������Bya9�7l��b��tnwOL��bq�{\�1�_D���kp�����=��8����6�ޞ5Ksg� j�7H�(Q���|��̑:<Wݰ�&$q4�Лf��}��d�kfU�{�{~�~ў�EmD1'�����
����ᓣ��<>P>�Q\�ds,�v:��o�s��l7擁6qw��ks_d����}s���A@��8ٹ:Gws�y<<���"Ђ�'3�D��lΛs5�z��ˋ�I
��!�a�7�NU#���⻜�s¨���������
���:֐�kT��j��{��f��em�
�#/C��(3���������m�ب�82S�GM�uw�r�m;z#;�8Й�aX��P�)�W}Q�v��YG��.{t��YUingU��7�=����N�6��%K���quٞ�^1sl��U�ws��2�X-��.��ʫ�5.R(P���u���n٣������!ƻ�δ��{�#�ފ,ķ4����0�x&�Dedb0�r.&^F],��i�7fZ�{���n%`���ޫ��u�b���Puv%�I�LWx��"����v�%OnmM��ީ�W���k�1�*��7F�t����R��m�LEZ�ػ�TV���.p�)�Mkʆn����Wڛ� �kv�ا�6�����A�v˂Gj�w�uw�S܌�d�%-1�i�Jܼ�UFjV�f�w��tD/c��.r�p�����5F��AC+�ћ�.OF^�q�ov���Bb\�bF�{�	�l8��3b�U�e x.�X�w�IިJ�l��8u��if��y��W��˯g,�mk���5�v�%�o���C�=_��^��Y�P����畽�s�`B��:2GN���/���z��M�#��̓��(CTw��cN�d)3A:��}����X� _NHK��X��5���H�^��}���t����5e�����k�D�:�r�ڶy�[�q��'��ź�n�Đͩ��N�y^(���+�\N2�;{��9t�D�.��xz�:>��;��~L��Dog�tP/"1bĲ��@�Rv��^�Q[����P>�q�kκd����f�3 �x�5n��m�2mR��؝�%��g�8�Bg�����#��k��ξ��?w�G���b���|3v}�n��_dt�_{1��CS��n��nk���:�n�QZ��K���`M��6���i���d���(���"{�?�_n���)���?�2��p��:�յ{w��d,m6������y�7q��+��?[5R��V\7�w�؜�G%Y��:�|�o�^�_�k*�Y�O"D(D���	�:�Z�3c�S���r����ws�ㆠ7�����Vvs}3������NV}��)�gn��U[+��Z@�m��{���o\��馳�gQ��|$�N�V��<"b�lį�M���K���BhM��E�΀>ǦM�4�/�{!DB�QZ���.D��0xFۓ��Ĵvm�2~���xu�3G>p~(��V���c,OΣ�"��7��.�e�<[��x	�:�,�'�V�6D�-r�c����:�8=]��W����R�3��r�ю�s&���l�i��]��m�76���`���/��k�X+vW���2c�����A�뜞ӳ����$@��TR
�A��uuhF��c��O�6J�7�"�b,��u	��(�ko�����[���u!�Yf��6�����ğ�U*����6#�_p�A�f���{�M���{Ѵ��[HE��<�gG��U�Q���π�B
~��������1�Q\A�W����S;a�WĔ����Z�0eM��
J��0$�&���;���t%Ė~_٣���C�ܳ�VE��Wek��D �=75�W�Z|k���i�1�X�=oWe��앷�W0�BwΉ�CR���o��^n�
��D�w�����i�b�%?{�����i��!_s=�Kx}��@I}��H�V @z3�e����fl=�-��^٠����O����x�Ud��;+|Y������(�(�r�B(����ʋaku��I�R��s����~y�Ѹ����sv��$�t&�|��zr�Ln�C�� ���G�BL�U��8���7�������xm3��a��3�!^ī�ǪQ�	<m�&*(�ڶX�vA6?�s�9�Yz2�o	̈́�CJM�����D�\IԓĦ��Y�B�~�c�Cy��$����{��b���] �c����9(8
Pp���;W�'�hVj�������ؾY|�-���(�k]�}����1ܰ�Dr��>��=��}hl��[J'���5�?, ��l��>^��~	�Y�b��3����N�q�j��f;d{�rC�9�ʣ�4�(�х^��p\�9V�ލ�	�����!�V_�Й_}�����3y����EP6�k�l� ���Z�v���v���{�̝v1�^|�ձ�/�xG۱|>�
I�J��zi�{��`���C��G������v����Q�R�/�f}��9��x-�+�݆�0"
�#|�L?��in&~������١m�N�t��b`��Xo��n#RV�2��b	�P���6��q7�9��l�1��vH�.��cm�턹9/D-�w�3��v�	�R��ٺ��l�=��*�������m��:z��vu�Y��̙��p����k�rA1䱷X+!�|�?���#n��أN)��'��γ�8��a��[���h��S��W��z!d���ǾJ��}Š��(��e)5��h�w���%�`�x\|����ۄ;v&V�.�?�h��=��}5{�o��u�n�(lBW���޹�|�g7�H����'-tdrF:��A�݄�Y
�RUj-�k�U���!o}s-��N��5�&E�����#�� ���}�a��"^P5��@�t[��l�ٱ'�.G��ggRU頤PQ�G�E"kjq!�64}��ž�8sn;���c��45}�������ꟶ>�O�X�����F���M��-�Eܲ�,��AN�5�?�~9�yI��4�1.��:��Uc"e-�H
-#�tpV6��RTeЬPa������ɮ��������������� �X��kb��1Z3�!�%kT՜�ޙ���щW�pL1SգZ�ݥ`F7�\��G��G��$���:p@��:߻���'g���5B�6�R[n�c��]����j�T������D7"+�r���N(���ğ�3�'���U+T�_[y�P�����IP�	�n{{:fwc�ѡ�v!�5�+�<����w�Y�w���}=�gd�T���V���%�b�}Y�����⏡6a)[�A�����n;�9�*&#�M�S���Ben�(�(��(}ad\D�������ˈ�����󵩡]�]�MH��fv?aht@���Ua�*`�-r�$���!�͉���o���'�?��m����_Q���jkduTh�i�#��lsu�1�Sڞ��7h��lje�4�z��$Ӭ��;ٟ]���]�����
����w�fc�w���	�I1'���NVho��M/�5f!)6�
��;�2�ul7����x�ɂ7�xr!��V�i��3ͬ��^��~�������WЪ��d��P��q�`����k��e�nm��?�O�m�8�(A�%A�PRHi Ԫ&%&��RJ*� �`�	fD����F!�hPh(�Ԃ8� F�R�R �e�L�"�Ң�B�R���H��� �T"$bD�DW�AW����E�Pn�*�jEw�P(�Q�
P�<bp� �R�P
D�
�
H��$bT"T(@���	� �.aD���V��1*A
���Ʌ?�s8,Be7�;��|(�$�%*���(+�ك����>Ӯ~>~߬�0�������������gf�?�!�#�����O�}��;~����>���|�������}������'���P�8����������!?���ؠ"�x�"� ��Ł�����������������~#���2�y���)�?� E ���0��̓�?@���\?�G��N�TJc������������DS���m������?����6"}�A�L��4�%0A@PDA0DBKEHA	!JA	��K�@A�$�,�00J�$�I��I�HA�I$0HL��@�#0@0J�B�J�@0H�"�"�
A"H�2�I$�)�0C@ALM�AA0A�I�@A0I�A�$AAA2��P1�P1�HP�!@S@PD(P4�2�
�P��J$�	2�B$J R�(P!!$R�@�D� D�@�%	�D�A@P@D�I0D(RPP4�
R�J4�P4�0%4� �P%(Ґ���"-
�*CH0@�2$B$�K(�@���#*��H0,,$,HB�$ @H$��@@��	 2� B�#���*H	!�2@̬�A(��	+(�@$H@$��K 2	)
�J�2��	�-#,�PU4�0S!THD��$�I)LIAA)!AKT4�@��%�(R,��ʒ4	A@�,�B@�BL�(�@�# ��,��C,@Ȥ,JH�IH��L A(�2D�2�I� �?��0�0��� HB0�$��H��H HAL���4�AR���	(H��� @�,�	
JB�
H�$#H���+	 �H�	)����	@�,�J�!��(��#"H��
�H�0�
$ H��*ʄ(@�"�A2�"��²�H�H�JB���,$*�2#(��(H2�(@�� ʰJ�@�	�A �J)"H�#",(J��)�(@�#"� H4*���
ʰ2���,��JȰ!B�(# B	@J��$�H�B@�@� A AL��BA)��BA	�$+@�$�HA0�0@A AA
A�2$���+)0�'N�A(A+����+�JA	� �K���,J��JH0J(Ф$���
A A+�0#2��0HAJ��A0D�AA3+L�0T�L̔��	4RLT��Ă�B44�APSPD�C-I!@,�P0@�"A A�0�0@A!*D0L�P�D�DAAT�3D4A�B����]Bg+��r���,�7����/� @:�~��~`|Ï�?�r0��c��=��>�����c�k��8�'-�!�@(O�0�������G���tA��C?����'��FD��v!�o���a��}���?��E�}���~��|����(�Id�H�����q�>���w��ld7�{�P,�� E �����e�F��k�~܆ð�`�"?�>O�z���C����@E �Ϭ=04ɯuQ@;��� plv[嗼�l"���������4h0�<�P0�NH��B�>_0���C�>"����k�|;��>Xg���t/��p;���?����?Y}�����z��"�]��#�{��  ����۱��������ڟ�c��Lx�?���	��d��������W��/���ք����Fr���Ǡ��P{�`Ê>�����8~�c������TC� ?�_��r<+��?n�>��|_���8��y!~�#�i���t �Y�:L�_���.��o�y���>Ǟ���?�B��`M��:�.�p�!O%�6