BZh91AY&SYҎ,S=N_�py����������aݟ�    @    �      (�   (         �=T	QD�R��*RI$��
�I"���PJT��RR�BJ�"U@B"P���
)J
ފ �R �� P HP(�$P((P ��   %UJE U( ���)J��@*��z$+�)#�[8�j���(d N����HtCA���JLtrh�r�	��J��(��x��W��j��<�'��� vf�0yuGf����p���m>������t��_{�t�|�����x���"�R�;��( ��K�|��W��xl'6�c�����<ڼ�Z�uQ<����g3T��:O��e>mJ�9k��]iP�T'�xkҙ�<m{ۉ�U *�� �|nO}wx�{�w/�Uk�;O��j���xl���U\MkJ��𪯉��n���H^���u�����:֕>���(�w�*I(�JB��"�� �T����o]5���4��C ��M�R�ۀ[����`' �T�������� J��R%*� ����>@�}��	����y���@�S��rA�����$�UI@�t!��
�
��à���o ��������� YT.ۀm��rCv ��آ����� 9RT�$P ��`�r ��"���� ���r !�]6���i݀IJ�!C��T��� ��R�P��R�Gd����;�j�W,�`�@hr �ݘ�uJ)XX�;� =B�U$� 

y� �� ʜ��{�@hy i� {�D�f�`@�l�;`=� �
��*A 	P   T�2R�@  �   0S�a%*�4` F� �`=��)@�`Mi� 	�0�6J�*�z��� ` bb ��*Tр0     % 5TL�4��ڦ�����i�h�F�����#������߿��������u������C?8� �q>@ �ڧ�

�7����~s����]$A�U����-ie?�@1P�A,�QTGR�y���}��
��?ȸ�L~;�?'�?�}�?\�	��;;��=��Y�������ŸG�
���q~�'�d�)� 	�X3_l#�1���+eDb��� ij�fHoY�51ԎK��4�KcG�ft9ҫ�����joq�@H�Ϯ�^1�rnU݉�kyta�c�l�Z{\���򽝽�-&(nH�ѤJ����=$���}z�q�o
�UEӅ���f�N��E�~�p�i�J�:�*^�=6�+��w;NLC��I]�b��(Xx�y뻺!�N�ѠF�!���(cY�x$��6�rU��6���l�XSC��"]H5*�T09����v4�M�L�Ύ�L�i������.�Y{�N%�a�F5(ތ��Ӌ��<���Cq�������ug8NT�D슷�g&
e�v�w!�;qת�p����S;u������+;[�]�-���"�����p>�������W{!���.v�ÄM�ȍ�]�5�h�2�ü�Kn�r�ь�9��P����<���fC�lrG����Y���q�`�v��^�lj�-}�4����SȨ��c�ٱjt'�p\T֏od�k8V�ae� 4,� �r�f���y�7+��m���t�:�7�1 U��n�<��Z�)�#`䵔�դ�u�����N�D6����#����V%�Ƅvޙ�jĞ���p6]܈��X�^k#em��D�뺒/Tp�X*8Z��+V
��cj�Y�wKG����)��+$��qhuH�K�3(	�;�ww���4v�4vk�&SϷF�b������洺�Ƹ��e�ݭk[%0��c�]�ӎ\����;9X暡�H�q���8��@x����A���5��; ����h�5T�oK��;.ι֮i���Sȹ�Oh���^��.�7��y#��Rq��v���4&�׸��Y+N�O�����Ђ��qP���BVYz�w�C�9q�/��b�
�{�sZ��N:�3����ø$$�i�q���>�Tdll`2�C/u�\��m,�Y�B)r���A�d`1$4��/`ު�:k���#$�
�-��(|�N���87E�;�=�)�����4�1&��]�#	ڃ��WFvr�8���.vE��]]�*=�����d*�� �;����;�����g>َ}�-�: gI]��@�����MX�$&8��R<��%��p����*b3#Nh�Y�C��f#��yg]�QU�05[�M���LƷBv��;�-��|a�kw�Q��4"�Fn�-�U���>Aǵ�׳A�
�\o�:Vtd��>�:92n��1�b�&ڷF���*�b���]�;x����r&��M6n��l��[�^�P��(��lQ��wO8�Θ��\�f��n7��L"�,�;w]�*�.`��6,zH�76X�/�/)��c[0� J��I�=���$rs��'#ۋ��n�l=t�2�͢�w)���)s��%�E��wb\�ؤюbS1d<���t}�4����L�f�ᔞ�GA7(�Ӆp{v.pX���q��̾e�J�=���*j/ێeQ�d����v�i�r�E�s��n��>���-��u#�@�4c���F�,DR؈��v���C1r�\���\믦���.ŜH�-���`z�n�y�GC�i�eED0v�5��CI�ܼ�75\EM��\��D|w-����?N!�H@�7�����grnہ2��|�D��Wg+l�{gG*�.֖]e�2��W��$��I�6�&(/,��op���ʛת�ge&u'd�Y��#�ю��bv�Sh#�x1�_.[�gv��n@���{r]ZF�ۅ(������$�;�9���͝Ւ���z{^ʙ�q�o�������o[y��A�]��у�w�����G�Zo%�Cx�z%��泍 ZMŔ9�Y�V�D]�\ɑG�ٌp�Uz���R�9�<dHa%��6<�D&Դ��K��PV���h%]�*5�3�q�R���^��@ŧ��:@�� A]��xqi!i�;�L�#4c`�[v����I�!��w�@y�"3��GZ�lg�^=���I<N*.�> ���&o4����ten*�x����N�݋����'�K�5��$D�(	Ӂu`b�"�Ƭ�P�s�p����H�L�W~f9a�ftK@�om�(z<�3�J-�)6��KX]��8'^�n!w����s;������E3=��e���֍Cp�mD��Ju<SL`�̕.]������v�Ph���Z{X����4��Uǎ
�(sXNسR�k�܋��^&�<(ZQ�4�;��{-X���=�5>;�"��Iq���(,���{�����tu�X����8>8×���K/@w�m�f�m��(h��{2rnhR�޹��=V]CN�'m��a�#M�o����8K�K9.���ooҹҹ�۹�Fn	9����^�dD��b���G'U��p�;�;�յ!F�Bt;��[@����ī��s��IJN^u�]�Ȁ����AZ���8rg��'̙9CT#VI�(�00��~�a�=ӝ��iF�� ��s]�i�S�M����uj9-غS�`��eivr����fC8��vXy�2�n2��MrKUä^�y���L���.!x���uŻq�9�,��ڛ��QЦ��؞�MZ��n�!�S	@���f����϶��ٗ�9ۜ�5Ƶ�p�>����R7A�L�.���B��\�2�<����l_��KYg�� �	ːp#�.�X���C�f<�k���!�D�[�_]k5��d�lX�����=�sA8��>�~�.]�7�a�ݜ OOb�<��;��n��gRC{��O���]���\귉�;��P�G�����j��8ae#�w![���{�wb7Lޣ�/{)J�sHG�\6�ꍼu��܉�Oqi��E��;�O�U��u�l%��5qԗN&#���9>�f��b܁ց;A��F��r������&ni*]޴�ԒQ�����1�FZR'�Hq$@��*���L���}�;N�˾db�Ğ�s�Ƃv��x�BN(��}0p����B��q�6ӝ�F�h��{0į�ǮQ�,b���%���P��B'Z�=ӻ�����Ż�����"*鋛��ΰZ�Rvn���4�s���	9�>�I�����`�9����0����;WP4��de�(��]EBJ	2 F`8wY�✸l�uCt�ZE*6d�#��T�5k�d<]�_jZ�V�'^̄�����hr�(�3K�8~]�i��y(D�r��Cݫ@f�ˑ˝a�oS;��C���uZuI[�`�3g^i]���^�]͉���t� �wB��P�d�8ɦ�v�7�q����➒��.e�
�6�����.m�[;Gl��@� � K�Y�B��1ecG����P�MO���ޝ%0;_č�E�Hw+C7��U��賕R�˨l���Y�d@G� �uvj&N��j7���U�͇��DV���y�֘�7���H�6G���"or�M��±�t�N�>rW�-8]x�E����� �� �*w5��!)�ʵ!"g?�wn�'UAj/6�ѡ-Ӹ�y�HG�v�H�7&+#����RX�f�k�7w�&���;@x��p�4-Y���'i�p�+����*�(���y��sfK�8���Nr�kS���q;�����:͹Cf���⒖����.��1�5�H?=��	�z!���ƙ��W��gp�������V�u������z	�O��娕��j���N���[�wf����s�Q�����x�D�"��d�P��i�B�W�J/�����(��/d�c��5ŻC�*0^i�ˠs{uۖ�7�`X����\�:����-�rFג�{&wG@y�n����Ӷ�0�/�=���ҟP�ӏY��\XBݠ7�+��bb}��p\���vi�DKۂV��`�o{����E�;�O�i�C���6F��w�2���w�����z�0��a�.�X�i�iʔ��)�p�Ő��n�qA��FY]�1,�]��N��ҥ��lWqx6���q]ݯ�y90�ݘ�pd�LD��78	μ��7��#$��-;�4��e�aV+&L8B�c��J��!�p)� ֐k^�5�G����!�t#���xH8�+9�kܛ^]���=]���K������V��ņHtԜ\�u�l���돚�p�-;�_i�{d� G��l�gM���AsX�*I1u�xg3'ŜK�rA��v�������ɠw`z�s+�q+N�12W��.��-YÙ��̓6c�o	˂��L� wq����"_a*�����s�s��Od�sŷ:C��-;�^w�a1]T��π�L�����>Y=�0t�Bs/$��y���=u%w[��K����®&z�+�׬�/gg+ۻ��-��tx7
�ڢɫ�����L�,}�k����Au<��N��d����C/y�''ae�
�c�4�VN��u�ps��.-���
�9�����IH3n��-�Q��-S�������n�hvs�7.�w4s�VY�ĭG�Ko=�2��Ȗ���7��Hf뮵��㓛@87pC��V���@W�gr��фA۰�Ӎ���$T�ONy��n���5ov��?��K=�����G0D�S�+�-�d��.�n�#q��dz-%:�a�̸�Wpb��8�uL]�v���H��JUf�W��}
�5�j�}:�Sn��_ͩvr�MvP�Wt��݄����V̜��!&�
C.V�ʄ̐�]_]7�g�.Gf�a�V�ڲv��Ȧ�m\��M�n��U�<�x�O��Gm�����O*V��ް�:؝���Tzb�&����ApN�qn폱���b�7�1Y�>t��l4�]�yR�I9tr�d���A��!W�Ń��{��{c��
R����5�ľ�nu%��x�׽�o.���H�.�ݺ�fj��'� r�l�2�����;�C���y���pbr���z�P�VB�f�����D{WeG�JWnܸI���z�1%�A�C	�ۥK�Lո���ױn��֙����)��:�R���f�T��a`�"́�E�Ғ���uh�\��]��:�6�Wn9-;ڞL�nA�꧞\p]y�dӗ�Y�85p{��l)L��V8ؔ�ga��Z[_d�,j�qιo1{F��\^m�5�m�w
���g�)ן 	|���FN{Ś��3xbթ�m���B�����3o(�����3;�n��h�uf�&h:a�^iS,�{�����B�r`a��eY7
s g9�(�)��
�ٍQ��� �X�#�i�a����t�����`B&e�&e���P��=[�a��F��»H���D�t�mf�#�n�oqx�ˤUAŴ-��8��:l�YW���FN�+�4�B�*��ӛ��Ռ+��=����L��n�3y��
�r;�W�`���8�)ɛ44`Iɚ\F��aK$�2-3b��7U�VrQ�)H��ջm��:S�\Bk˂�7r�x�}�,�X6'�����OL�铢���0Cs�P;p��{t胏%�٣8. �9z�Tuv�� �'2FWH��[�)su�A�n�I�ԳM;���Y1��mf�:.�t�ewU>-�X<�.rN.йC���wf[1<bs�4�� 2��dh��-��N��U�f�b�A���֌�ب��.=r�5r����O��w��wks�*�Ѐ�Ǥs�o-��Ftf�d{�:w�X�i�ɡ:�g,*�y�����JU����N�(rH4��N�Y �<1ɸ����;�9����j�_�������N��O��;�{F(�8����eT-�������?D4�X�~��c@
��wm���;����ˎ�D-tN����iJb�K�^̩l�X��y�G@-��SFQf���B�A��mK�i�r�j��(�a�e��V�Q�t02����K#.�	n&�C5u�2�)�ƹ��Š�vm��)�����[!6��l#��3�P�ZWktln!P"�%�]U�:ֳD�FP���Ùh9�f5.�"�,���1m�rCq��K�9��jGAԲ���itդDG�Lf;)v"�-�N���Mm��\]4��,���/j9�SK��&�ũ��` �h���Z�tZ٦�fVa)v%�c�G�F`e[	��Z�cTfR���ԺTv5� �a�����w3hE�a�t6ve�q����ep�jde4��r������]���ea�+�����k�e&e�A,�m�띱���8�h���2��Q�FS�t������FηY��Q,��mh-���kl+��	VJ�ȸ�:(�s�� ����	b.3�Ė��bB�6Յ�;���UD�2�Y�B�Vm*�T�Ql����ccv�[��\,Ε���i��Zd��i�M	R��d�fd%Ŭ�B�F�Z�[�De�@��c��F���jK[�X�K	rD{��kCM���_3�&$�4���[i�����m�-5��)0%Թ�i%��a�5�5�ƕW:
$]wR]�,p�7.�-"���a�\��4���eU�`
;Wa��,n-I���h�mҺ]'.q�:�!\���>n��EYH�>Q��\�p��9�s%K�a��h��t�a4n��Kn����K�Pf\�D٢�M�%�kmͫA;LF �4(iMQ,,3�I��*�Q���BH����m.Gp�`��.�uq��X����r�\;�X̓b�t�a�7Q%�.f#,��H������x�a3o�z�˸���/y��<m��z�r�x��kc�@�С�`Mb����^�d�J�Ʋ�Ɔ�`h��-Һ32ւ@&��`B;C�Y���.��e%�V8{Z(�)m��&�Xl�B1
M�k���j�6�6Xk�2-"�RQ�kír�@�ilT��f�Z����)�(��˪�s\�f2��]����0l^y�n6�j����-5�2m�nV�2�\�J]+�Ibk��3tȱ5��u1����z˥���Hqg)YM0m��k�e�\�uʓcY�xH�r!,7#'�Ûh��k��dZ�U�9�k�0��&j��(���nՐ�B�
h�6M6�F;Q�!@�b�V��K� �Yp��Fb��,�\h�36��#XӪEm����v-�A�k�v�U@0��*F;#4��mv�2%��{R�J������Y2��LT�z�0��.GBX�a*�R�Ļ�,�������[���d6T�յS�aiMΕ�QfiH�jX�R�꘹`i�9u,sZ�1](Ҫhe֪�,��Ўc0�)�ݘ��!b��Z�X�nB�F�UBQߏ��]��띛1
��(	 �rݱn�KSAe��و'�1/����JD��(˵�n�`Ҭ�4.Ơ9أ��8�ĸ�����
R�[1�\��".��[�j����X����vmʎ@�ͺ��U���[BՏwj��4�4��@	Rn��VZ���hh�# h�-28���ɫFU�m�:��J�+R.�jV���utv�q�0�B�2�M6���M�
p�E��B�5�M�Dӭ�`���]�\m�i�ƫ�LX8ֹf�U����RʹV�J�@�R�6�,��F�������_<��F�+V��IX�n��5��@�-4��Y�l%H�x1	l� ]­Ys^�ŪFө6�%����K5�i��`�h)[��(��I�0:��'f�f�r&�:ˑ�SL.�4�c	v*D*�f&\�K6T��*�&KeJ�e!134��Jd��2�� %�L@�	��nƹ� e4օ��܌ۺk6ȁ4v]�n1]YP��;i�-�aAd�B��6��|m(��kF5��kTke3p�6f]Tl��z4Ά��:�lb��J	b�mf��kX&HAi6Я7*ۈ������c ��n�a�Q��X�ҷu������`�����@4�VM�x���{R��R"8�;X��Z��Xjfٗp�%���J�Xj*��`]b>Y焻����`Y��\��������4�n"�貛�l@S]K��1r`&�+k[/�x������m2�

 X�ds*7�
��i��1�[-A��pf%�hWLf
�4V��۶�Xǫ,�X<����S��$���S7q����Mv# �@��u/n�����!qad3�z�4%���6��T˥G\K��rFƨ��gJ�YPZ�5��p��k��݅2�&�GL[F�v��F&+�H�t�A͑����5��v���1.����8p���:�.�-�&	JFWYa32�0¬��
��%��R�ڶ�I�ʶ����l��9�n��V� 1lk/V��4Ҁ���uJ9�Cm��� �3Eq���f7]h0���h��f��L���I����DJͦ٘-�m 6��Uuv	eZ.v���=�(]�G.�f@{P&f����͌ZEp��E�u�ƶ5PP��\�������2�|��b���5Qt	�;b��	hL�
@��+3k����MJ�k�;@.��y��I]h6[P����<n^)* !�9�R�,��o�U!�r��y��:�:�my%�%����Pe%�	hmra��HC�E�d�9V����F7:�`�m.�KL[f`�m{$,Ԇ]�*����YtYDs���WמP��h.��f� ��Z�% �-9��S^F5T���m�� K��mn�kX�R7MU�ؗ1��.,�C����L������a��k;�eO��qm��vN��-�� ���3f��Yn�]g�
�șK�0Yl"ʅ������Xc�,�Xv���r��!.��m�H��ZGV�+9���q��y�SJ� Ҍ�[u��#���!���K6�� �D�-���:�%��5 �hsH��B�A��k���)e9iM�\9�H����.��h�0&�iu\�Yb���UD��{,hBZ��`4�4�vڸƬ1	t���̭�foX�d�Ac�ͬ5�-�D��l͈f��ћU4y�aŔ���ZVia���{v.%b��t���MD�d���FST҄k�]��SlǫB�f�3	�`�i�Q�X����;X琺]���fl�K	�bf�v��Q�6a�u@�F]X�R�FV�����A��Y�t���7��\h
K���h�B�:���Է�8Qp�h��h�M���j�:/;�BT�]ۇHa�����0�b�N�&�RV�Zxƣ�]V$$��B!�]��J�c��77��C^U�P��32]�p����W�#J�iJ&�,��i�R�6�f��j�b=di%	rkm�W7 �F.�-���_<O��f(���Kll�])-0�i6d���B��c��+&�[tt��|�4Dbq@�ԥ55��q0ҭ�����`Mj�f�QVm����E��ʥ{F-F̜��.�Z��������]�:ڳ1͆�:�C7t��M*��i����-�LڳIt\)@�q�4���րl�7v�f��Hr�6iV��5MF����BP��nn{9X����кe�ECU,�L
X]o�̻C#��o,NH2�1e!KfYk�cgS����tk�M���Y�A֍j��F 4�LڭYp�jl��$�j�	�����Mk�0��v�n�	G�CH�v�K���5�&��X�IKp��Y���h�]�YJMt"V�' �]t�V��L-RP4�iV���Ү�K����0�iCD ����0��A�`SA�W^ͦ���X6���K64��t��0�����tv��������*3��5Q�۲����ƛSM@���=�M+��2�iR�e�+.p13�C�	�@#o6�.aR�m�T�=^W�6�<X�C6��;k���L��$L,X�6s&nn��U��1v�`�Ut�؋� �x8�]B��p�5�%[�v!.���1Ý�,2�s���Z��n�7����,�E���ͣ(j��;&�0����j�אd�6,��v�5��.3tɚ�s���m�V0q��7�[�9��m�\3q`�@�+Ś%t�f5v���J�z�ذ�I�����K,�cf.�Zr��&�Q"SVvѷA��d#
���l��+]���T��X���)ζ�j����F�،��[���m:=G&�\���ζSA�]-�)ML�d�b��q�Qq�a�%����^1sR1k6aX����b��!��X�R
��8�F�.E�F�v�n��6G[�Ѧ��a�Xbm��q\����̂U.S&�Ѭ�"�Ck�G ��v��K��ݼ̑��ATG���.�
9��v�DC�7̟�/�/���k�U��o�'���u��X��(h��|�6�Y�u6�bn;mڻ�pF��4��������m�iN�f����*��;�Yk�o��id{TDj�_1�����lrvu?x�_T&v�'��5dS�r��;����~9F�L�T5�I2|4��S�/U�~~�ZY�����3q�zb�sd.n�=pm�'w`96����wxzx#r3��ϧC�3�n�OF�+&I��z[�'`�3w�pg�>�o���y���w��g2��n�|��|��.��9L �x�wՍ<�݌mg�23�;M�ثĲow��%�A��Ww%����]���w������k�����a������xn{���Htgr��D۴O�������K��w�!��!�js���S�����=q��<���8��]>�!<���O�Z�v=�7��
�z5Ux��Nqf������dVꞒ½�(�����T%"����<"�������w\�_\ߤ�[����6�A���9���8 �����PL�q-�r(���X�R�o��ս��>j�?xX{�NK�H�2�y(ԂsO�'����w��_��3�Oh�w�q�O�~p�qa����"�͞s��
7��r�F���s������p�%��s��5?N��Jy*f�X�5
��n���D��������1�b�HT+��+I�L�ԯmN��\�ٻtUN��Q�{����aB�E�1�>Ҽ�b~��ݛo{͡�=1��G�>��0�ن���ݸ����2z�*3�<���<&��<�=�^���yһ�aC���>��С%���xf�}<}R~=��Y�J���=B>�g������v(�E��� r���3�)�-���y���Oyw����g{�ˆ��f�#�I����K���{ǳ�l��c�&x	뾳���
��L�r���N�1�eLlY�p�m�w��~�:0�>�&5�R��w(�Y?%�F8T4^��w��'T��0�HK��р�s��M�C�OO���쩘W`P(�K<��=��~�D���l�"V9D�+���m�o\����=�݈%����ؑ��d��K7�A�-@��mޜ���wy�ۣ�D��-;٠E�{D��14 ����.��on�0㯼���������>f���͘z)jکʜ�Q*�e�&7St�lf��h����H�4����w�?:K6!�tT]lλ������:&0l�UXA�J�ܫ�h�xq�f���m�ٳ�[��f���ȫ��}�]�twv:=��V�ai��QltitZ���w��=�q���7�����/rp�ꆷ�k(���}��y��N�ı}+�kNs����FȘ%�v\�{��V=ȭ�𐝧��/q�3DW7�x�.�2|��N�����sx՞��<�f�q���ub�KE����mb���:�w;"�ڄƳ��g��}�l25<E�m/vW/����:��<F����@���Ow|KuF��[~���#l��T�U���PR��g۹b�z<&͑d���7#҇�)Ys���pPl����o�ݧ�f��x�$��z�a����y��{+�ۂ�h��'Q��ǖ��/<7A��D��c��k���ܶBHr��\��ؓ�#�[���j�������*��=��y�I<��ٗ�ԋ�{k=��G^pcs���x{�7�N����j6���9�����-p]�0o��r��g��i��}��}�vp�+^�����ZR�l[z��Sz��z�s�hE	��J$�ZRsjq�[��L�ݻ��A;�-�����.��:E��-��x�٣&�f�"n�y�.$���wV64��u�9;��{�r�@��'���d���z2�U�G�����v;�PR㈜�M����Uw�K�1���l����qvx��8���Wd�����{��?ygdl�i�|��Z�R����ڼ}^S���E�{�Ո���/�|�q{�
�oze�8�����\~�W����i��ޚ�ܫ)w��]]���N8x(϶�ű&�t�rŜ՛��,�(�[��s�u���܂+�p��GN6���4鱗`<@�o�����7e���� �44@,<��ՋR���y8�m[���Xw!�b�t�ف�3&�ݢ��op,:$V�Ƚ�~�k=g[1�0�h>������KW�eY訴b�����uNs���@�@{@��G�=�9�iiM������<�6A-0��Ta����2����١�:�D,é����	lϩ�֎������ڪ�0VL��=���~�A�������8�\��ǧ7N���L��rW����:^�	�vm�d�M��o��b��W�]��(�.��N�^�+[%ڙǋF��ߥ��_>n"�^�������_�ܼy"��4�k��٪l �j��uZ��Z� |����Q�zr�9�!�7��xlS�v{,�S��I���]��B���g���v2\�tvξ����y�$kMys���[���)\6�r��Ƿ�(|��Ek>?#��=8���5 �����柰���靹Վ�g
t��x戽���-׎JϨ9�E�{��&<�g�+K�Gi��8�>i^��Ɏ�1��դq�ー�O�k��T����/H�q�iQ��j��4�˲Ml�o+��7����:{�3�x���{4h}��u�i����p��Y���_���ǻ��1�z1|��sh�Ƚ�Jb��=㏩y�4J��D$���׊�g�ۗ�t80�����h�Gô� \��|D~& a��Gc���B"�y��Nz�!�.e�w��;�����&=�/C)~����§f�Pn�t���/g�c�&���ub݈�����k�f��r`����3����Ľ���J���V`c)n�پ����8�JG�ĶN��>.���߻���� �X0��Qt���mk�������*	���v��'�.j�\e)A�i���͡)�&���_�����4�Y�]��\��w^�>�4�
�4!���t�x<|ր���|�]<�����b)���E���3욚�6��gi�7�����kdS��3�}�����v�0zv����.�<賳����~�짯LX)N�Q�x��u�Sm%���.�ꓙ#��-N���׼�j}2nw���P��1��y��=+g�wL=h������ۺ��
1��3�g���	�{�]���=��c�����c���K�
'k!DǾ>a�P��Rj)�mV�'u��{�@�,F�!�[ѩE҇��kf��f�ב{=7�m5�y���ʙ�k>���r�p�vw�w�{�� {��ڽa����m���>��inPAܶ���zg�����M5{�ZE����m��쯖���zS�v�>�d���wU.��d�*��zM��a+"fnX�#'EcB�pBݠy�h����W�u\0-��p��ξ�Yy!���o<:�$J����X6�S�؝���*�������}�m���6����`]�x"NZcMͅ'|(Ó�u���P&ߺE���̚�p��=���q��'���˯ ܻiح�ֳ���x�=N�M�@g4��C}B�MEn{��M�:�i�P������ŕ�K�!4�����3�4BP6��ة��N���&�u*<s��{f��n�n��Y�Y�5k�"�~�Pw���Y7Y���7�E�UŽ�l=�F=wI����	s�ꐟ�B{Ww�d��t`�xێ�1��l�A�����g��ZE x`�N��m\�Xb@wVv��SCL�;ی;g�9��F�Zܵ��LUf1!}���Л�4I�o=��'[=�O�2�t^�����yU��wt��(Ȧ�'�ޙ!@o�<Y�^�$:4�/pI�A�;��];�&�j����7T������T�'r(}�z�
����h�tՋê,����;a�i����{'Yw�=��^�K���G�<~_ww\*�(,����}�z#iE+��"J�L*ӂ�j4�ٜ|{ۢ� \�'����V{����.�kY��ܘB�b�×y�o��J��+�*Vvļ.j�~kY;����, ݲ�����M��檽���D�^t�zu`�6HR
��2cro޷}_4x/'��>��n�Ҳ)qox�P����H�Bw�U���xu�q=-�>Y��c/�`z���gY;M�<�F��nn�"�M򕰰nhU�u晃}�:{����w���OD��\������ER��n�f?r,+���Pey���������֗z����F�BABvD-�wL��d�(2�S�-��@�,���9�[��/.��3G�9�{�������z�
�ry����.�{�6BG�5j<t��<w�g���e����<��Oi�����=���6Y
��(5s��K*��OME�!����O�S�n��n�B�TӋ����.{����wx�t��?O��=�����F�#��5}�'��n��|L����.^v��A��M��~%�ݗ��f�p�<�:���!��u�þ�;����'��[,���sP�P���;zb��(��1�!�����y�Y������?��M杔,�������k���6�eE�`�s�[�3��<�n����3sz�s��Pɏ7*�Ƣy��X��Fǃ�r�U�[w�����\8:sg}9v�|�N4y����ڍ�'§��i����F�t����<'P^n/ d�b��X7���9s�=,�nn@�M�鷙~��ɶ��{�� m*��B�fA�You\AX�X�P�yL5Qz��V���r��OUF�ۍVF:�����k���e�M�Ʋ�?$E8���>�|� �����DL��<�/���]�|c��jo�戮��s�o.�nNd���!�/1`f�E���L��9��)�D�g&�`ܪP�&�s3�dﻒ��r�Q4����xwm=3����+b���6��9���榡�&����;Ru
q�a�x�Q3�#�od�D]��N�, �ؙ�;�5ލ����N��m�ɛ��ݏ#���jUU�4�E4��Ӱ�e��N�ys�����r����zN.{�8�K��n_r�y��Uㇽ�\&f����N�p��4�yv����Y؂�wP�������D�آ=��%��u{p�q0D�{f4�,բ�G�:N�,��a���C�y�4H�	���&bΦ|E�!ޱ^�b���Kѷ:��nm\OqT�M8�DhK)Ti�+lx��i�����>�|��Z��n�%�g#Ƀ�w:0�kE�-�r�1g��(^N�o���;����^n{�zu�
�=��,z��|�{�9�K~<`����3����^�`������{�JF[�[w/2/�!!�7��t�o�ᶾͻ3Λ�t��f��Ύg|s1�-G���d��(����0�}�V�tX�frJ����Y�g��Jwx1��1Ρ�{����ɴ���Σ��E�^OG���v�ʒ>{��{�Mƀ�����g�}t����l/�4��G�Cm!|=��^�8zk�^�ho{��^�:� �'Ժz�*{����Ҳ��x��m/	g�4޳�h'L�;�-���&��T�h`b�
o'�֊_|��ss~�����	���Dn�4���m�ѱ�[N����I%�w����&�'��;BG������ө���� �緯<�V�[޸K(�و����Aж헙CF*�ӵ���:��3���w���=��}3<p1!������^	�p��w���)���｢oC�I��_w�#����F9���y���[�/oa�#�Og_,?u��?-K{�RS�<Vc{^���^��=뻆��0[v!�>XFY-��ίn�>���[�
����G��������X${'yT�p�/}ؕ�����񼅐�]�ݙپU����n��/?m����"�d�b�פ>못pR���g<�]N��]N9u�^��6�h�*6�J�XI*��d������5�7�����j,�����W�gh�������{;�[N��]��y�'�r�uN���6�f޽�1���3&E�{�-Cnj����A�����}�L���\��GsUMq���h��Z|3٭z��uGG���@'P�1�!wIK$J�� "�/�������U��vA�������>$��B{S�;w�����P�6\LÉDUv�Tˋ2�J�JJ�t%s(=�	Qu*���c�kTil�b�e�V]��V,7E��j�ݮťe���LFPȩ#e�KL�X����m[dZ�wXШƍ�Ļ5љٴ�m�n�\�)�e�3,C�M���HITŌ�qtk-t�tPkH+��+3����V3�)�5vy��,���V���L�L�.z�bj	f%�K�f�b�.�M�t*������W��4p�M5a`��Е�v�&���"�"ЮnM�4Efs��� ��Ĩ��;l���X.�0L46v����s ذ��ń��X�\uj�b���͉�kp���ڔK ��I]f��l�k����M+*�iQ0���n�E�5���-E�Z�Z�\�K��Y�A�٢-e�G,]��68�̴
��[r膘ҁ���
2�E�Ņ���lѩr��+��d������ɨ�u��1� lE��D� ;�V�1�Tqu��[�r�\ZhW]k���tl�RU�jGk1u�"�Ť%Zs
مZш��j2�RgGbR��J��\��.�XU�=EؗRG�Z�%�i��4M�`�\�v��r�i���4f�u�L1eC5�7	6DVh��-��j#��khJ�nv�
Sb3V�,o.�r܈�J�(Ka[-��è��� k[�������fvњ&�SZ��NF��q,S��ױ«7iG���!mf��(ҥ���R��ZlK	e*�
Rp�6�nZ�#���F3�4&����\��C�49��m�f�\n�,a]vE�o���)v��#l�*B�3Y�0�4D6R���+Fƨ�16���f9�7\B�2d��"F�m�-G0��ɜQYEh���#�XZ�T�Yl��������ʞ��+'F��;�W�6L�Ȉ˺�H�Hh�st2vd�p�zߒP�W۫�Y�f�uߨ�Ϋ��g:�R<{�F@�h���ƓI�RrH��V�~�-�Y�R����q�������|���7���=�tg���k���٫pg�M��l�E�ab���ˣR�}s��L�*�v���ّ��������ݔbM[ͨ.*w⪽^k#Z{��IZ}*��^9�G�lc�=Wf���g��zqEĭ�U)��j˯h�ve�sO��<����9+\Yt�٘?o<��`�CRTA��sj`�,u�59PD��TT(:qŃ�����c3f�a�)]U;vcq����Y8�m'ϓ�0�d+H�kڳV�b�3|�7W���c��dx���j����d!�R1�M*�b/TڡI�БQC(���٣,��MD�4�a]�����Mx�&�X`h�@���X?e՛�;���`�_8��=��կL�dn  �wU�����t���|�7��kZ�����t��<�jvQ��)���'r7 �
���1��U(D\L�Ĥ]{����Y��yg�|~}_��!H��Vݵ�J��4��B����v����JR݊�5���v��#m�ܱ;iu���6⫕���	.U��z�͚i��cS�eЫ
��]`��]�DF�lڪ���5��Y	�f���]j·�l؀B)�u���1-U�=lZ7B�!+�v�ik8��HMpX��WV9��c�zY@���P���ӻw���F�e�uh �m����!V�Q��+�D��.X�twh�Ka�(��_��][��P�K�t%0� �8,1SH��W|>�ov&eݡSJ�:�p�	�Ҵ%�L�p[,�&i
Ef�q�B�}������#��SK�QPJ�4ڊu� �;�\��ޡN�j�1<>
/7�j	�脂l�I��lK�̑;K���빴�bfQ��4��lE�A�[!�qG�tЄ1iY��j�.����l�5�(��e�� ��o)�J�W��i\f���6���U-{82Xl�	�ẚK2'�#X�n�,�Ek�ʊ�g����'���6~3�4��	�W���~�_�z
�%��3��{G���l^�^���I��7}���z�צ�{�$[D��l@AF�hT���N�j�5���ڎ%��MCi���ޡN�d����L�����x���3`���#E,�{>�]���o)�J��ک���-��n���p<:�QH�sE��sg�/x�4_zdq\gP�K��<�!D��I0�� �d2���ں3(b*GMpY�`F��LL�Z�Rܱ5Ն�����9���E7������w��oy�!��A�4��Ю�|*�F��t���H�mW}�[|�s	�	�
�n�m��<��s��~�ޙ������ݾ��2&ȣӋj�cc�����:����Lm��Cַ.�V&�6���ÆƯnr<�}�� $��$��L�9�B�����8-6�4��\ y��T�oUM+����>�wK��
"�i�E�u4�dL���\gP�J�p�J���=* �1��bRe��Yf!#�(����kuF8ll�,j�)3��Y�)���T���|վ}�UK�tRb)4a4Zb�+�����j��ު�W�+� M���%@B6���s��ik݊� g:�9F�t��Ƹ%B.P�l�6)W}��7z�idoP�K7hUTz�Vqrޡ9�OEB�����NDUĺS�ͷ��V�n9���9�J��vL��Tpn�`o�rX�ѱ	!α@f>1#�D�{54��$�&jqSH�ȗ+�yZnmf��J*�j�;��-�6����K.����h�m�]f��` M3kLk4�h��&ȣ���G������ס{�3K^�w���;2%�ֳ[1.��l�Ҽ]B���sz�idoP�KwhW�og`��*M�M����T��| ��i�����*Y�%E��jN��}�Žb�.�3=��.}�Sk#bI�*!�Np�0j�jk�fw��ɤ��2��Nv�#���=F��X����3Y�B7������'%="co��VlΉ��K5�M��ʼ���`�(��y�L]wZJ4�
��L�;=j��]H���@U��&��f��̠:ΡY�]Ql�������6�6�@���M{D1�"%�j�#eI+����l1��L5��2��ф�-�0�B⒋kMmR��L3j0�3ml��$ưl��:���[R�nx�.JB ��Ȥ���&0X66�Ҭ#�YbaQ�Ք~��a- ��R�Km,��=y5�)���A3�������̭��\M+ms��T!*ل�Z�aGg�ω����ƭؙ�Xǀ��5}�4���QIC"!6)RW�=����fاK{�L���� �̒ %�Bh81&c��L��x^�������n��cN�L'
�G�=�wH�uT�כU�|gu��X�sL��i���M,�:iR��6*�\fЧK;hUR�Ψ1&	�"Hlp��8�[M��.�j��x"���6D��\�%�w6��EU#��*i���uo�OT�x�taBL$�8�J�6�l���.tH�����
r�Dm���^U,�G��f�BɁ.�V6*62���gƞ�4�I��2xg|Ǉ������Ds6�ik͊}:ӂффц���sg�M-�:iw��ln�L����[���(AH6`�[5� �;��=誤w6�Mw��b施fr(�f!3J�W�.W}�bݭ�UH��z���;�~S�]�E�D94b��؁��5���jK.�x��U�ڭ݂˱L±j�ߞ����
�W�)��S��ݲ�b\���aM	1�gm
� �G�v3a��x4|&��j�.��*��TR��B�c#�Ng*��o*.����T�o?~���� 6���{�.���y��i�ú�ө�}�'�)���,�TJe�bD@$��|�E*Y�B���vK%��E&�����E�#��*if-�J��s�6�v�p�H'�m��ک�x��R��b���.V;Ȫ��$f���66Xe���6��S#���/b�mZU�B��U��hahj���1v��χ����)R�S��"�uw�}uo5uD��i*�1
j������Z�bff�sk:� �����b""bTZ��U�f8|-���"f3�c#B0� ���GoPs���n�Ȕ,E�4��m�M��܃����&x�#=���Eq����{-:1�6�T��|{O30�<�YsJ�klDlvuqϏ��1�An�UDj�'D&�����ڪ�9�B�#6�ur�����s�j	�3v�nc�c��6S`v��c�©�V��0ef��m	��n ��_����[<>R�ު�\�@�`��"�13y�B9yA�f-�U�vD���Z��l(I��-5U��&2�j�c;�T�f�qqB�8-MMi�9��1oR��$���<>x���L��q�ջ���lux��7�1�qIݎa�3��m�U�i�j�{#�hki����D���lD�E)z�qk�k2���D냱Y����xY�eÒ�K�DMQ��\�Q���L���]5��ZK0iP�:��ڸ@���"�F��A �a���	���eإv���0֪��Lh:5ɫ����Ɩ"�R�[X�m��궖f5�$i�[��G�n�!��ͤ�I8�i)���,*Z�G]��\ۄU�զ���t6�дH��#�1a
Xs�|Ք�--	hu-���xAc�u�st�D(kS:4�˂���1����,�Sa��L.��ZP�LlY7��&�i{W�
��"f1f�%�)�ӆۊ�;�#��M,ŽJ��H�{�\>�Z�zO5S	�Luo~m�;���>�w�Z#�<L�?���p��%�J��:;�S��7��<>3:^f���D ReBs'2߾�r��[ԫN�q��6�\$��`�e�i�`��l8&��j�ɢM�T�F*�4ٗ%�wq��bb�fdVd� TtwC;��!#0�	�
m��gN'��U<�g��I����J��a�d����:�C"E7g�H�[)���#\��Ӂ�~��I_vb�B0�@� 1�5ozD��ٓV������%�Q	�p�L�wH��[�=��R;�A�f-�Uhdi�B�D$��|�;��;WLL]����ݡS� �䂄�,�*�sdL�}��z�����ʓ�������a�Q_�	i��zf��!2�6���u�pX�uQf��`�W�s��̑'�v;��^7]�Â%&�Ai��:�|�ݩ=��$��|>;�I��m�E�s1˺&c/&g�� %�|1ݙ�Ri��}v���97��0.Ƈd��ؖ�����j`�����۞���i��񱊄��������:݁z�S�z�2sԦ�1�$�r
�:G\�EZ���߹��߯��ܘ}������o���8�Gߥ1us�S�>�<���0���L���L�a-	�I�b����_!�l����]���!;�ו������ng�5��xC�k���I���c�.��3ʇw;�5�7'wO?g�{l�Ӆ-�+����� �|��a[��U��U���v�9�|M?�@1]��w�Kٹ��DG��*d�J`��יu��d����d���ӌ��q��y�]���<����8:�����o��(���S~�T�͂����t�! �:a[��\����{�l��碗p���Ww��3����ܩ��<�>����t�j����)�[tj́��Мp��wbj���1�r:�ŜK�m���g�՛cbT�ܱsF���Fg�z���s�f��G�;c���C�P��,�)�d���ۍ�"6�B�ۈ(�ΜFTe5�/�޵��w��P�qw��w/�?zޜ�E�9?y�g���Ϟ���L�p�_*�V/-^�J�l�n8�FƇ��%�:3V��k��L�"�=�)4{|\�� [�E�ݸo�A��מ@���+���+:�с-7=h��9r�/�� {��
��膠2���4�p�8�52Mْ��m�e\DA��(�C�5��WI2Ļ���x$+�×ʋ0T������1s���t��]�ia��2�2F�����o�z��x���`�fomE���wgM��V��'L7	J�A9
�����û}���ϻp�j��5�0�/�4�>����}� ��]ɢ3�:�Zf�ܕV�\n�m&wJ�}�������4K��9�n�;�q;��]X+h8����Y�{y9��d�A3�`����3f���C��}ƿl�y摜u�';� s!d�T��BD��D��jV9��ta��\�1VX�=ܕM؂Lٔ�Ý6\���N4!oJ�omӾ��
�!��c�Vo��&�b�*�r��
�"uB�I�Q#%HD�b���sy-W�R�*�N�g=�4��t�(��[pL,�Ѻ<p��A�d���2o�t��>O�(�j@���+�W��N:n�[����77eC=/�G�Csplb�I�f�^r�^�ac��8#42f�țG��t��j���4e�%�9;��=���Ω?6�Ww�ŧ D�n��as�U�!�����'��~/BR�@�[l����f����czɸ����&���ǃu��l�I�L�܋??����Mo#x�'{W3����u�^�Vja�O�F����!0���ß����3�MGhRU{U2�-���k+���}�^�c{����ߥ}�k3m�B�T�jiFgf�7	)�,Àʺv3��`�5&n��z9Ñ'k52��x���������wF
;�����Y7Cq=�b׫b������LL��C?~��|  a�����e1B��j棨j$�{�.��wn��<���jݰ(9���{:{;����)��#�c�ɸ�P�OZ�S.�������O�F����A2a0b��?WY;ڬ���Z̎��>�=0���:w��K��QP�(�uO�ͧ�u��7�2e:y{�vXx�a��u��{d��ڦ���.�`S9�u_��9�ߟ>fx@JIN��)�l��������O�~��`$��jJE����O��id�,s����s��b��pf>t��~ωYm3�bն���V�i�l�[��*�z��V�lv���-й5���N�F�0���ms��f:����GZ�������wS�|o��M��Gks�;�I�s��R31�O{ՃQ�^v�Yu���x������8aBpQ�����������Z(A�}ZȒ�V �M�*8%�I�ට�'��/=ޟ����z�C:�;�5wՄ�^QV'�U�lֵ�|e���0$���=����|�~�������c�+�:�N�SuS'�=�Y�1+�C}�@��)��s�����<~閃���u�c��b�XS�"�0j��6�D0B�b�˄c��[n�Ў�l,9�M��m1�dV�RU�GW6Ǝ&f�TjL@s��ڷ[l�@
X�f�CDhB)x���1Hִ�)I�3�х�4�(q��&�wi�Sэ����mF1�Vh���l��nf�KfM�^ʮAQnu�YY�]Vi.��9�ڳ`��H����+�v�~B~��R�ҀJ��|� ���2�K,��QHi�4����]�1�L㰚���(�9b9������������M۝�Sy���>
M�;������־-0Z�����5��a�j.�^���U^��ι��<�w�z�`š|I{����LE�=�˨';�`iH���`��{XLŮ�><`��1{�Z�˨�!�0$����L�[�� uR;�W��#���y��l�I�M��|	����0�{�&�o��ֽ��`I
 �g��˓L;F%\�����d�Fle��!�l
����,Pe�ՙ���{:~_��tIW��_�ɑ� Eo?��{sBRa�E�� O���<�^8�Q�?�,詃4-�꭭pH��Z#�^���r��.���[���܃��3�fe�cm��yGk����}��0��I�b�w��_�w�и�CP�&79����������zp�h)��-��n!�� j�I��5ݳ��y���QQBfpT?
?��I��}���[ؕj�aI�<��S��/lLb1����V[��3c6��lV�
)��V�[�v[�48pچɆ����^{ޟ���o6>���<�}GỾ	?}�������l��D_u��ұm�C5m�e1[��~�<���_63�nG����`	?���ᛛ}�"/{<c^Z�a�w5����<�<��ɫ�����?y�hO��N{��{�~��G�?כq���GNמϰ���I�A�#�b�I%�KoW0�Wmq$3�X��v��{�bּ�/�5JY9~�e1|�V]A9�cR��7�� f';�Z�Z`ŋ��%�/��3��{.��wָ��."fڪ�b/E����b��10^������H9�ÜJU6��uf�5.�g�����10�P-|cN���9C{ｐ5��P�t~�����D|;�A��@���>��@�"�S|�N�1yڭշ��gAJ�6~Df�R�$�be�	ˮ�����O��BR��u�mk��b9��^���a�$��X��c�b�}U�.��<�Y]F����e1B麶=�s>�^T��7���O���Ò�yx�q��,��w{Q��S�9�Q���Oh�F��'�"��9�T*����p�~ �����@d�����=��N�<`���5O;��N��wru>��t޿?�ބݹU�Q�^v��.��4��Ϫؘ��4��smL�`Z�4n�l�u����iWT�(�]����.ٗ#���gR~o�~��;�Ӽ�j:��{'�JP����}��#hw^a�X)�.�����=�}���}U�.��<�Y]F����e)R.c��e�I�bؒ���MGQy��L��h��0���&#���*�=����>��(���l¬�>�� ^<�y]D�U��N��Z �2>����-��-�n!O�Q���J�M{��M�1{�uo�����A�^��'G���r�M���X���y8L�3�Ʊ5���s
2�j
ߛ\'c��`轙jN�F�8�����@�`Ě�b̎���&�.��2���-Mu�ڼ!Ib�A�<�u�I�85�%Z��y�/ڵ...-�ڦmz`��n6p���Kb��K��j�r�b%�k��Ճ(�u��k �[,�٫���WM3)l���Rc�>]�D�/��)e!E�	��v�M-��Ch}��-� ��b��$�9���-O7�ʮ,�]�J�cZ����+���2���͋��lLZ�~wp��V���*m�M{��~~{Z��Ϧ]E�}�g����[}�����C��l�)~G�}�+��|�[��/ꬦ#���}�Q� ����>��V�j��yގ���}���;�=�m��u��b)����`�o��}�'�?!���͇� �s�(Є1c�Yy�q*�FGQw�g�.����asC��oj_1y�Zז�1����';|��o��'{�l˸���j�k)�j7���h�3�����F�,����q���&Y��Yn�h�GU.t��D����pl��h\�Df��g�?�����&����;씌A9Ǒ;�C~G��͒`F�	0b"b~���=�S��&�˕�ok���F�W�l��
������z����<:����Y��S5vXZ/��Ԙ{ٴ�&wxw��t�I%�\CT� B�-@2�a��{˸f;��֌��^��p�b�!������6�IÈ�j~E��;{���G�?�&����}�/"n���YL�S�E�L(�!�YP��dI��>��`�w��kU2�&�x���P�(�I�~���~Bz;����w�G�+h�&�x����l˸���,B�U���7C��V]�1�O{�0j:�xR�g��Y�GJ�f�rU�@-&�K���z�gZ���Q��뇙�a��j�w����~�zz'���;컆�����`�j8��{�������G�~�Ce�$���M��H���}컔]G�*�fGQ/v�S.�n���a)X��X�X/�0ч�ӟ��?Y�w)I��#w6��d	���qˡ=�v�B�t5�p��5弻e����eH�����E1�E�Q��X�N]<!dK[|����-���x������z��,���\�.;qHK�� !	H�Z6�{�L�Q�={�w�q�/���K�4[ls<���w��N�'��n�^D�/��P�ow��S1�(Rt�>?��w_������.�Y�z��^6�{YL�Q����f�/!��%Uh����I���˸���B�����<������%L��%�R�γ/Q��jU+T�ӣw�F��n|��=��/�ߟr���w�Ƀ1�Ký�vd�b�"a���~E���B�!Ph4�%7�p�w�����Cp�9��L���^5U�&����;컅(AMǑ+>�P�D!"�K��X�g�d#�w{YL�R
�8�=����#��U�Z�������u�fu\U<�gOd�$�;��[�Y~DGoz~���ğ� ���qw��[R&���c�tdڡ��N�A���TμV��ެ�lc�h��w��;�^��1��;�C	ٰ��#),���ϯW�_=^�r+�tI�" K��ĦъW5��j�����w���ď��	�(Gͳ��m��H��"��O�Gq�`	U[0�;�xs���wp]�U1�Ѿ>��

f (�(8�&ѣ�����t�ل ��an����9���sp�8�ߚ�y޾L��^�;�.�n����J ��!�b�.��'��ы^�/|bIs��Q�K�|��2�PQ�1��P�osՇP�u��L9��"tN�>��_��2�nY�{:{&:��Z�f����˸b��J�كq��Df��g�?!�lI����8�������/�V�1�Nv�0f7�xo���wp�@�z���5Ý��}զ�V�g��D�gO�>z��w��)!��s/"r�Uk	�j7���a�~�����3��*�ͥF�U�H]Vm��O��.��d�t:&����;۞~����;}��K��]��k�7��}a�v'��;��o��^f�$x�Kj��X�3��6yEmd��Z��3�>���U�ʭ"�h������vG���5���y�8 �A�ͷà�m)���w��"��|�[�J���Q,��n ���=:7L�*v�õڷ�s���Bg/��Q���hxzN�p�2���j^D4om���s��,�pAM����f;�74�ꙺ<�m�|�Dy^_3���z{��9]yVE�g��kX��2ߺ�9@�]NN���o��dվ��i�	}�*>U�D��o�Lr�<�ᾜ�e�6&�ȼ[y��ڭ�Y�Ū�=�
٬�������f#���\���s�6A��ݣf*�$Йo��)����ɣ��r栕V0�B�*��#{��.ּ�M�GTиY�t��F�l�0dD�2w��vqu2�Q���Y�A&jE*�W[j��WZ�!p.*`ݫ[����c2J{��5bʃ���/���Y������R۸�)ϗ�z�a�Ūb��6��vk'�{�:�7ī
+,S������*U��-�A���S09K�{���ε�c0��nJ0�E#�M^��s��MFB/qLͪ�S1�;z&^I\���~g��niBE���]w�7�u_�ry����;l����_�ƅd�.��Q�L�MGo`���G뺽�g�>�&��&�6�sX`�u�HJSdo�v�P��;P��au(n�c�Z�E5�Gi�KS,H�m�ֱ��"�i<+��l�3[.�젱�)���lCd���3�s�%��ch���Zpl�&��D��)n���(�YV����zƮ��%�0�U�in�NӋ�����f�D#D���`
�++`[�]U��YX&F�	�,����
f�X�$�sM�.����mq56�p@amt�r���9��W1	����h�2U.�Ⱦ_-��L��[a5�Z28�A݃	�z�6i�1�)H3V[�- C�m4KT�`��`⺒� L���充�0���L�;M(����L��F��a��&e�Rd�(�{.V��+[�h�RG2�`¬�i�С.	[3�,��<�3h�U6!s���+�kʯX=e1��tq^�`L�4�jC�[h�!1Q�-��Y���k|+���%1�m�3��14.˴�-)U�yk-H��3�m�tk,�ԫn5j]GD&Gh����xЂG3l���
C�뮺V�惣�����5)J�Jb����m6Z:�V�����Yb�� L�3�.1J���� ]������a�!�=I;� �#�M�3��P��[Z�sJ�SsI]l[c³ 2�m�UлW�1Rd5��Filթ��������Qkc���s��$��-R6��1�6��Gx9��֚6XQe��$�p���P���{j�V�Hs����3+m���թ��:�Ŷ
):�#m�6ݣ�$��4)I���%XiKv/k�r`\��ȳ�]��],5�6]LM	�eE�m%���ȗV�����b���X��lh�#-����1�*	j�B��Y�tm�]��L���8J 0+�ꈬ����uSn����</Knd[,g*���s�І�C5ݽaS�6��8N���Vy�4�@�Y��8���dǹ*�kBޙ���%y�=�8�o�3p�i]'&��3�i��h�BRn�R�.��`��q�N�G*d<���t�(�W�y��Q�#c���Li�+:d� hh����܎�įn���҈;��B�>s���G��0���[3��s��g5l	f�	��SL�UW�����wfws�wC��ۧO���{��SF�F����7̕�7���p�7$Z��*>i�F�9�wS%�z����<�����)�\��D� ��/�v�(+t:�9g�Pc!&���{Z�'�.8���䱳I�&����h�P�a�i��,!Eg�|�|��b�>;N�m��J��'a��5�1���F}#���,@b˯���Ɛ��9��r�t�{�,�8b��[�GԦ������:���B)OE�GG� '��(%d�v�����t���h�܍�-��D��.Lꩰɸ�6��n:�!���Q�q�����J��ͧE��!��� `��tN�8�qQ�c��&�Z�����%��jv��<t�T)��cra�H���/C�m6���.�+�<�4uq�^Kbg-��F�R3�
r5LK�R�Hf�n�-���5��.*�S.R]5�,�v%�����i��{VR�U6-GH�ł$5[�u��Dnl�I�3,�ã)*��V�FӝA`Q��LV�0�nz�%��>=�fQ�;.��l�-eH�al�Zm1vcm��|HI �����%�h&D��bI�W*�JP���^�cn�z�v��ʧ<e�+��ѣ(Ҩ 1�ܥ�n�������(l�ʳ�Q�K½�ٗq7��ﵔ�5�}ǽ��NC1�J�уQ�K±^��(��h�N~������� ?dY���èf:���&��/�.�x�a���(5���I1	�����G�Fs�e�1������R�C�j�e�����?�G�Gs�-����Fc�F�w�уQ�KÝ�e�M��w����(E1{5YC����� K��D��G�#�E�u�����G�`�V�;��x[��&����|�3�Ͼ���������da�YvX(�1�2�j�J�Xꛊ�-�z��x(O!�¬�	߁xڽZ�����{��1����)����#7ޱ?Y A��o�ME��iBr ����¢��Rbۊ�GM��G��UCˬn^��f8S�����vs��pXR	1�y��ڪP�e���>o���z��ϟ~��t0h�"bD�����bD(���3%�آIӴ��o�����߫�yQ�w�2��x����n�!^�Z���&�iÈ��!����z�U+��~���~����w�����
L8m4�!�J��#��{]��UU+��v�� �����]��W�%�	�a1we��XCQ����U�p�w���d�q��{[2��xҵFj�w�r�Z�%��\]G��Z��!lM�)6�`�R�Xű���$�C�H_6l��r>�,���~�g�~�>�{FGPo��ْ��� ��Uk�E��c�����- Y~�>�w�2jR$@u�\2��x�լ����=��($$F#�=�}a�$�ؑG�#�G�ޱ?YY������������ҟߢ�]S�	����ӳQz! �b�"�24��r�<��
�;I��M^v+s[۳�E��
������K��Su���Y,!G�~�H�i':�r�B	�р�K�I	�2f3&���wU�w&�I�*�al�Xu�Pjޭ5��=��b���-k൤�1�pi
-��V�cho��7�������XhрN䟿�~��N�t��*��Umw����;w13�w~wFJ�`���ywp�y�k�j7�	]�W�[�1y�H��F����f�Ѡd��j���uҵ�����'�,B��m�7 a��}��(�Dos�ٗpw����R1w��o�D����.��h�MZLH����;����P��1����5×�VCp�w����D7����C	��s�������SQ~DF�0*�#���7��=�V����|~_���n��.w��'��I�Ø�VC��w�Z0j:�xo�צ]���j*���}�l1A^�9��צ�^**�ݵFj�L4�(��q{"�OX�طnc.�e&[�ĩ뮞��Pn��T��S�8��Y	�F�d�
F���$# �1a$$H��%�B$�=������}k0� �PY-�D����7�H����4�A}�W���^=�k�j7���{ Y~�>� p�M�b!�pPPC�zŖ��fIVlX��h:,�j��v�g��$�.n&1ic��q�Ý�T˸;���{XCQ�-�{,wGpyn�FMG0o�A�)m@0؟����~��`xCp�q_�Y�1��уQ��|��2�� NC�}��.`��%�%�k[�Q�-��P�uv�td�s<�PLC��p��;��n����5w�����Z�iW׳ý���I�>���3�����j�]��/{���� DQ���"O�G���(Q0��F(��7�{�ٓpw�R���G0�nF.��"O�G��A�?Q"4j����3+fnA7�G�{�;8��mʎ�U�#6w�5��#������t2˸�y�L	ޱ�18椼�	
6뉎j�c��\��\BŹ��L���� �ݭ`[�#��k�]6�l�f��D�/h�Ԅ�r�	�r�M�ͥ�$��l�f,E&.�e�6���V]0��l�E��3���
�.E�-���_B��<�P�&�&��k�q�]G�lK4�1rk�pk2B���t�ZY���%sB%M�޶��YwW.'��		#z렲���L��2,I(`���[�is<����M�R6�����5@Y�.�ZX\���Γ���0��[naU�S��/p�{_�uF�y�������� iP�Pq=�V��w��z4\��c%���Әj7���{!�B� 5A���5A�9��L���^>����"�Y~dn�	�ڏ��b�,�?Y�գ&��7�{�l˸��P��c{�#�"�Ȍ]�HD����7�2����%�cMGP(B(!�s��Ų��x�V�:��x[��P�u
B!�zċ?I"=�`�����DD&��d;��nw������=U��3D*�FGPo���˸;��K"��OE����4R���X� ��.5Ֆ�@�E���6�q-w�;�M|�y�B��k���=��ov��c�;�;�&��7�{�ْ��r!�۾�dsF��k%�V��r��p' Y~�>��Q]�f�a�)uO�ݵ�7%���HɃ�N��t d������b1�Ԭ��=ӭ�`꣣OgH�/�u��z��Jf$,�R�����&�T�'�\Ȕ$�$ B�A�C�2��^�i5F�y��HTGp1���\�MZLH����#��b~�>��-��k+�BU���U��3���(������D&�ٟ�����P���wF�{U��5���5 ��B#xUz�eBѪ�x�`���JG̊?��(�?}���{FD-��j�x���D�v'��'����٧�e�[�6�ĺ-G!)i��bµk���v�4�!<�t<�xmh�I�1|d9G�{�֌�� �罳.�����k%@ 5���U��3���w�D4�.,@i�~�>D^N���M��������j����<���&�HD�C�慨/{^�!{�D6'�#�!�{�#�"�ȋY� YE��U������P���|yO#a��~2��7�������Bh��ߗ')�2'�t�<�,EX�ʎ�3љ��c��>�w����|b֑�1��HB31�r,9�I�sF Ɋ��0���!��G��!�?Q"/������G�y;2Lb�ėŭldsC���{U��5��Z2j8�x{��̻��RP��oz�}$Q��w�����e�a�ɝ�=�h����
@N�^�wp�}�k�j7����Cp�w��z[E����̭�j�I�F���u�T.��a�U�R�S�	�0(�p�i��ċ?2>D{}�wp�m��Y�F����d(Rr#��A�?Q";����"baCs.�����`(n�!nW�!�j;�}zѝGo��ٗp���b=��Y�@L�Nf�F��sk��Ux�b�n�^A�/��P�os��~A���B������gu������xn8�xz�[2��x۝��9��b��������k�'��2gdVpCY�u+Or�V�"ޛ��v�S���7�rŸ��)��e��ELUg� ����I����,RQjaA%&,�m�W�>z���|#�Ҽ����a�ؑG�#�FgWwp���U����z����>�]BE�"<�'��B�3$�2�f���*d�Q�m.`6�5�V�"���w@�i���LD����ѽ���G�E��7�p}�h�BCqý�����ؽ�G�hl���#�"���3����.��V̚�Z�V���Z6�}���$��z:{��˾Z3:����OD�����b����e��/{��O��oHE�G�B\�mC0�j8�@�\C��ᗐw���k!�j7���{!�f;�*�f�po
�yx2a��ۇ������~��c�"�yK�+Ր�5G��h֌A�;��d�d}d#����g�۟�^���z#s6���]�$�R�je���)�<�	�:��"5T]�����;k��5		�����tӝ��K�V@4DB�]��m�Q��Z]Ka���	e�X*R*�Rl��A5���y�U���i�a�	)M�:,�k���QJ�� �K��m���\��-S�0lm����tW[(Ui]j�]���vP$��=���LƌfeH�v��n]�vd��e�4�J�$�����n�1rځSQq�c�Dr�t�	�� N�J7v�nnc���LIFF��snX�d:@'�`%����uf��&�	f��:���4�6{2�f_���恊h:�o'f���|=��3������7�9�l��(�!��V�:��xz�Ucb��ik�1k�!�j;����2jR��C���pw���k#�j7���{!�}�	�=�N��>�6�+Yc���:�xw�[2��x���R� ��#=ސ0�?Yo/P�G�GȎy��pabIk��e��.��,
b7��f'-ꬦ���{ܘ3 �0�9�{fPQ~�t�2@��DH��G�o�����1A�j�d�B��z�e���;�dsF�o]��ykʾ-b��lP��X2Qt�P�X,#�k�0Ħ�(���/��KMf"-�D����z�U,��d}d(���
F ���r�Zެ�c�b���m0\6$Q���#{z�ޫ�2�I&/e)�ڵ2`�6�ь�����y������8����ĽǓ{S}�#6sq\U�wUâ�ro�6�ˉ���$�I�@(�P��["��aY66����FJe`�I��S��~~{�����W��wo{�0j4�pq{^$�bCl(LH����g�g/$5C�A�}[2n!hz�Z2��h��ǽ	r��1{�1���r��ɸf!�Od�������2���b�~��J��q!�d80�w��G�#��5A��`#��p���x�ٸ��ज़��'�#��|��{�Npj��|<��e�����Dheb]u2V��Q{T(��M��F��	���bF��7�~�U��Z 3�B������P=�9�V���Z���T�k_�%�&�c|��&����}송����3k}�F����~J�4L8��}$Q���DQwz�� G�D[�����'j�k�9�7.�8�<��K��0{�W�l�Ϫ�]���*vdK�ĩy�O3&ӎ�mf��_�i��U�����I��`�%�[8+�^���_ �n���"��ȍ����R��ܵ�ug�h�7Ϻ�wn��5�N:q�N�Ŷ-V0�ϧ�Ao��Ɂ]�Nt����>��k~�)o�=��+�Y��M#�w�˓7w�R�Ox��`x�'���<x:g�9�}鰗����z�([����^��������;+_=���`Cz+I��n��t��G^�zyM��>���Q��8<fg�+(����޽s�kn>[V���\T�,yV��s���X��}̽nk�B�9�S�]�w���0
D޾y��|����y'�zr�|fѠ�obi@�6ED��]�v�LϝM˩-j���>y1��[7oW�K+���0��W�6�%��]:q�
�e]��08m�=7��{ڼ�����h��zVQ"w���,��k�{Ot/$�s�n���b��jʘB�f�-�����^E�a�}M>��>�9�/g���f�ES`'�^��x��<�I؅������2Pj�=_�����}���_�}V q�W��&	K����{����!�N*4���c�;/.]��8V,�"�-�h�Z�'�e$]���I�s�$�0��	V�&.힧�n�r��j?���|�RiM�^�ޘ`u�f�>��B�$X63ze�jԗyP��t���F���=fDZ����]߮����-B�jٿ7��X��e�r0��cG�n,��M�N��P
����2;M���t��!�(�ڴ�3�J@ټ�v;�� �����$���f"��A�A��3V ��s�����o	듲��t���#�=���R��eዏ�����7�}��;r8��ֱ��w6v���u|�#�Ws����sS<��.�7�`
9��h�:��ĵ|�H�W[�k�`��	W�.�5��I�CH�~�=���S-c��S�������D�I�D�z�����g�C�(�s�$����~L' ��;���rOKI�a=�b]*��٬g�#R/r�G@R�!�2�a/��]�|�����^�]l��������>�v�u����Ghd�
3�T3[Զ!X�!)�P�AFf sбp�ӳD��4xN7�}B�a�f���~:�P�~Zǲ�C;���A��[�!��|�����������8�1�t��M�:F�AS?C�mh�vPr�L�:��Vhɧ�z�.�	��1`��Q8j��v�`�M��P��77��4 ^����0�^�[0<{���=v[�ܴm*�ch��&�,�0��k����ʊf$M6�բ��5B~���g!��'�W�B؂Æ���CP�~��}�����h����XqC��k��Cp�B�ڽ�V��ۇH��F��	�
"������𪏮7�@�$���bO��pcL�Yn6���^��Zn��tlh�u�64�m*+�5q�]��ωX��ng��l�ׯy�7�{���)�w�2��h���D=�h����"���Mx��(�oPbO�A��5���>1�j���N(p'5Q��&c76�w������sg{��5xw6KA����Zb��|~n��*�u�'/*�w3h�����:���+a��s��R⢃�A}�H-j�)F�sYj�e(������]]]�9DOd}*vWnw6�Ͻ��z��	���a$`�F-�cbM$�E�A��Ѡ���BcV%?uo_=�z��r�e�0a���7�.}��}����M�v􉘻ݡG���<�a(}B�T�fYFᴎV����u�QW�]��G1��-�pf�{�2{3z�{zG�����ޙ��JB�	���圼�� ����q����Z> �=�
��I�[b�=�"f^Kﾏ�U��M�}�oHbHFcJ� ��6��p @���z�f߻송��w�ѓP
*7�w�09��w��ϱ	r��Z�CQ7nײ�b�A=�h������?DA�wP�H���3>Ռv���˴�<ff0#�ؗ�}�w�婜׷}�۸�GX��;���o")*��tU���ܛٸ�9Q�\���v	�^��$�b��5��[tfԖ�Z��ah�b*I�)
+e�l���$��f��`��0m�f�u�d�˛�`�6����.�l
ؖ�\��L��ۓ��4����J8�������)�nMb,aumW1R�����"�`�8%�e��#���3��.	,Fj���m�`�ak���8$�' v4h1���&��(�ÔX��4RUSQcرR)a5$X�Л����^<'��c������-R�.��Kn*������.�\̿���r�B��|Xd�ې(�?��P�G�-�0�ah[[��*!���k�D�c�eAE�$[r(���� x��-{�'w��s�뵓Q�*�pc��Ӂb~���y��~nw�C0�ȌA{�0j!hs������/||�qc�$WL �;�=_}���-]�d7D;ڭ5�;����Ӻc��ߌ�=�}e�-�-��C1��0f!i�b��̡�Z>�9�bNo��j�x
�U�Wmy|pvM,V���s�أ���C�٫�������I�R�Ce6��,��w�O�T-o�����s��@�r�{�$������a���p��?nj~"*���E�d��M׫z�d��{����W��w���l/��G�۟�/��x��{t��Y�1��݈���v.u}��䱠��{�V
`lY(JH�h��P�1�E�#Q�cQF���mtI�޲9���{&����h�P$��G�҂��,CEDD����� Q�{ܘ3�Db(��k�Z�����$�7P�l��paC�ZrQ������`�R�Փ+&�ہ�yH"��{��g�x{͒�i�P�0ؑG�"��5J(�{����;��!�j!�W�d�R��U�kT���|L_��є�R���Zf�u���qCG��,���W{�;��|w�Ch�`�g��;���4�:y�~~y;o�����j�{�Cp�{��W��ɫ�-|K[#�j$�;솥!�C��ٓQB�U�(j��� EQ�G�}�ȡ�LB��P܁D3��!�?U�����v~7��&T�z�ffQZ�+3IܭWy{%�b�f��t�. D7�8MUq�{��\:u��>M[������5jpŐH�		�0��Lh�֓̤*+Bwm�#Ih�*5��Ѥ���Ih#&�b�\�QF�Ub���!��'�s7d
"��j'67R�&1�&�Ұ�+�[2��hەXC15���C<,T=�k����Iy�
j�U<�=�����xO	>I!n��n�s�Z2j!h{�ϦP�,w�;����6��K��y*�13�t�Jep���q-��8�N����<H�!��k���q9��d5D;��������=�)B����a��9�f�Lb��-10Z��Cp�w���dԤ"�`���L���^6�V�9��xo���� s#��苒�D���"��GȌ�W�� ����`u)	���}YCQ�>�^�"�̏����n!�l9wt�1��y�Q9��d5D;zC@���@S�w�+���N����6v��k8vt����È�;�c]_u*uSPr�v��[��r��l�e������h�l3*)*JR����,��,T_ms%�(1��Q�h�k*Ch1�$Ba��w52��h��H.�$ك�}$Q������� 8���W�ņ�V�e���=�ds'��>������qW[n��d�V%Y�(-fBV%��%�\�jf 9��o]$���X�`�d9G�kգ��7���ze������7�����n���ݫ��yCm��i�~d|�gW��� ����mڭ�sF��qU��1��}�Yﳡ$���>���ذp�sk����p�j�XCQ�-�w��P�b��|�bE��"=������G�}((=��kܽa�B�C��Vy�nz�`�u��=�L���K+���]�Q�;U�y�Z�B��r�G�#��(�$7���ku2�<�j���5�|ǽ�x��=�w��VdȝjV�7RcN��Y��w��ܐ=���Ѯ���g"����=r������Z�ȩ�ρ����o>�]|�&/ā��G@Ϋ�A�&�����m�F�a.r=�[��\C��d�.2����QLK-�Ѕ0�ᚉ�Kq��82�K�.�[��X��(�6�6��I�A|�l�K+p�Z,����.��hݍ�S:\�Av�Q!/T*�W46�:�k(m2v��W���^E�5�,v���M�Dq,�B�2�?I8:@�X��L	��*)@�m���6&	�ͤ�
"� �C��@�!	!/�ys�M�cJ*@,��Q�TQ��v�m���wa��3c&���O����l�a0ZbE����~�>�}�k�j7����/��r�$�F}蝉������h�M+��󽓽�=�`("���s���n��׫FGPo���˸PH$yG��W!jlB�I~DFwz@�(�d|y�hɨ�P� �=��L���^=�����"���TM������g��e�[0n;�xs���w�������R�W�=��r���$���l����|[2j:�xw�ײ��BP�V�:�hoݪ�n&���Ʉ�B��'}���-rf�u�++TS[CMcm��ɣu�;E����_]���x�s�e������oO~�8Ĵ7�������&JF*��#���?YY��1>d(l�	��9I~D^����;�u#vTJ�J'��ݣ��y��յw�f�[�v�^�X���͙L\�d�8�u3�*_��v�����߿�&!#ɡ��&��QX�d�2�%�$�K}��E4� ��k�Pj����7�9�T˸;���{XB$���䟟~yw�Zh��-j�'�j;�;�ѓQ�þ�2�%	NC�V�:��xsت�n��߽�z�q�X��^���̚��R�;ڮyp�j�XCQ�-�w��Q�(�۽�,�D|��#��8jlO�G�K������5�V*=���!��z�`�u��=�wp�h����2P͸����ke���-j��.�l\e4�B�6�w !̘EL(	&���}$Y���p�ws�ѓQ������Cd}d3�guH�H��#5�B�%CD�Cp�w�����M��;ڮwp�j�XCQ�-�w������Tzi����������ѹ�#�9W({�u��qX�9��{�0�Un�f�pn��sp���_Fg�4È�K���K%:����@r�P��k��u=�g|ݧu�g�d"20�#$E�3CI%��s	#3D�	Bk!24��!�`P1�f����u_��Cp�w��s1�ø�{qu�i�T��w�w��u�'rw߿}��F�+Ր�5���5Ġ#�#���G�B?.=((=��HBX29��xn��d7�p)]X@�˛���罳.���{�����}��f\���Rj�.p1��"1F]2��b[E�ir�x��Ԓt�|<�m[�cs䟐�y��zѓQ����:��^6�;��$QCq�9Ud7�po���/��-L4Ċ?I"3;�O�|�| 9F����5�ܯVCp�w���d��g@��I�9'�?~o�5�%�J¸˸;��j�k#�j7���{!�f�9��棘7�9�l˸����v�/
4�n܏��>�� B�w�"��=��FMGos�0����V�����~�.":�3��*Wg+�S����������c.Ԋ�zmZ��N��:'A��&mb���[�fg+�n�"sj��e�b2�1�0���b�BR �@�#�Z��?_^�K�x]��nM��0܁dI���:B1z ��{�3�<��UZ����m���Od�w�wޒ8��O�ˌ�6���!�Q�DΚ�cp�)�kF#IY��7��<�����6Qpd�q��FA�/w��G0�oߵ촬��yޭ5A�=��T��">MD5������ G�Y~d[���n���׭5A�=��èP$��߿���ϝ���0��w��v'��U��3��}���@�\C��ᗄ}d#���c�"�ȋ�\!�L��������5жG��lɸ��]��:��^6�;��a�x��1꬇!����"(JdC)�P[BE�����'�#�^P$F����7�ܯV]�Q�Nj�(���c�/�G	�_E����B�R�`�T*�$�N��l��^�s������{�S���i7š�1�F�Qj�7hsOk��bhs��完���<�����n�o��۶�Rj�8�aU�":3��:lu!�orooo�~�4�E�gk{�Wu�&��{9B�7g�fTŦf/��s$D>��V�gq�U.1Re���#�sc�NXƃ�Ur��H�4xl���yc-Я�o1=�Ӧ���nZ�����J}����9=t-��U�j��f��T%�z��&z�ʻ���i���`�t��7]��R��q�s�nE=l�9�$��)��t������"�1�n�&-�A�Edk� ��I�z�fS���)�W��ʉE�d��E�۝;r4*���U����V����A�N1*Gl-E������D`�H����j�I���-���ώ�������b���k�IOuu�ǭ��ݍH��-�Y9�k!1Q�ڣufn��m����}��Y��k�d�e7��Å6��z{{�ܫ�P��a��f����i���G��	�;qhܨ��3���$N[q��x�+)[:��>)Fr>ۿv��.�L�]�U�^�������{;6��̽i�M��7�2͎`H��#g�O��XN.�_{�U{��e�o2^Xf�v��	�f/MC�u�����l��\�Z���H�@�cj�gi�ML�θ��0(ӭŻ9]Bʢ*�.�3�5�.,�� �*+l5��RRK�)�@B1�٪孙��Kb���k�	I�ؐ%�fá3`\������e�`uP�lR�.,����	@;Z%�]��!��R6^5xL)#Mt�6�,�a�,��J���L�����Q���Mɇ�qR�� ��P��[�.��j�b@i)(ڸkc��u�i�n�%F�\�i��ś�f�]MK�r�KW�4���j�)�e���h���eæE��[��l�jv�i��v/R�:4��,���� e�6��E7e�3�qv2�k]�r�q\Z]`�b$�Dn,�ev�J��*0�v(��1+e�f=� Ŗ^ƩYeЛAE��&�^����%l�j6��pGm�j��cfh�g��.�fkB�X��cZ�[�!�ڥCBj�V`���JZK�d�rB2�W$iL;J�X��Z���h1л%W�sf�2D�lNĳvP(��6���%L-�h�8���U+e�]k�t�q+N�@Ɓ)t��T�e���-��j��f�$�3��Ɉa!��@e��f1��s��q�����Ѥ��Kn��Ζ1H��Mt+
	��Bê��D�!r�pX9&][Us+�f!��u�!Z��.y�kK�M�ZM0Ͳ��di�4�`�ح��B��Mf�cvZJ��b;]����=J�E%��"��l���v�f��#P#��ѩ���bmbZ��.�S	��m�4%aJ�c����h,�����Ns2�T%Ҫ�)Wi�n�M���+��+e����h.�[�m�9�X/j�4\E�l��e��fh��ڶ�
�m.���f��`��Q���nl�E�L4�}{W�|f�Il��6̎�6w�J�G���L��J�5�t���;ThaЋ�����)��u&\lNV�ٍ l�R#%<��r�����Q����؏*,�'�Ǉ�t*�0te�WA-B���Æ8I困��%����;f�|�d	
}���,���� ��,��Y�4LCAa��%w�m�C�Un��Y�|E~e֒�z��|�{�
c׹ݼ�����3���#En�LnNiaeg��4�͎�Ѻ�b�)!�	�{r(A�i��<����s�t�8� Z�sq"ό���8�0�E��DKЁ�$�Qfd��zh#�����V ����,>��Uk�~�Zx�ƽ�a%�7��h�����D)Ab
�b�����c�a�2/�ߍ-{u���@�
H��`��Ɓ�G��+&d�!�.-�7�EnB���w�&���w�^M�z~`55��g S#��]�3��!�;�������Mc �#0����N0���K���Y"�5�F�9�t�pG�/'n�arǹ�:>�h�ji`��u��k��ҟ/ �nh�T;�'|��<����Y��[����,���ks�B�����C��HP�;��1���Υ���M�fq6&.��!�3V(���@��1��+]S[f��t")�H��G-]��*�2�T�І��9i6h����ř)cm��X��<Ev����IQ{8Z˥�M�mk�S�B���.���MayTв���f+̶���K��U�a�b���ipX\�ZZ9�N�Fk�k���l�k�,ό8�8 � I�Ҍ �)1&fB$&�B@ȱf��$I,]z�שC�b����H&�m� ��ن�l�y�mASLﾋ%ɉa4`������ћ�$}$To߾�Cp�w�����;��w�������G���B��l�Q#�"��w�������r��Ȇ�}G�}��̚� ��a�B�y�d}'��{9'��>���Q�[����ޭ5A�7�{f]ġ`��#�i��?"#�z@�(�d|���C�n �ؾ�� Rqw�0��x����9��xn���gP�b=�`�w��>��6e�n�)s<�gOd�~���xO�� ��;켆�ȝ��FMG/�7�O����<�������J\����D�K�Ik���\Sd�<WD��ɼچ+���O)�������'9�5D��{^��Fd~��$���uɄ1	8�6l��W�OݸA�����t�]�с�ǌ��$����(��ޭٲ��UC(Olf��F�h�ųqG�I2s�dn��z���=~_4P3&K1�Pc���kIH�!�6�4g�_Y}��~~{���B?FgT��� +[�W��>��O��&?�P�L�����񻵻3> S=�Օkyz�Lm��P��7u�>�ڽZ��=U�s���F���Us^-j�b�i6�o�/�z��> ��B&;��wcw�f<>�p���i�؀��i�FZ5�W)jՍl������ڮ�]7��͔b����|�wzD�]�uݽ��W©��뺵�O��0�L�ة�ݽb���`������z�mn�
� W���>1���*C��ݮ陔v�n�w4�;�d�>B���'^��㰌��U\K�_9����GpceM�[�'�."���0�����[@�p�������7Ѹ{em�z��I�tlE�К���5m2�I4�э����̡SK�}b��l�D>��pۀ�����<{�VM��P��������|u:�}���l��0
n��P���=���]ު�W�w6��Åz��Q�Hw%����j��H1�	������2�R ��i_S�ɖ��[0����-�W�ݕ�.e�����G��*if�4�y��A�b�����#귑�T�n�
�^��&���>�f^��m�Q
*ioz�ޡS���~�{]��ꩥ���y�m(d�iݻ��0;�b��wkvfe�Wj�|�U �4 �-y!��-'[�^I�4��{BTMt�/�GQ��b��f�Om�.w�K�eQų�0YF���q�b0XѴQX��Ih؋zk�b��e<��������C�n �1J�gu��^�����3k5uR���*�w���>r�����4��e�-����&��=l+ZE���T�t��ut"� R;~m���e���W0�����^|=)��4�N���گ||�;z�U,��b���Ͼ����bh�$���Z�^�J�gu�� 3�����]T�-ǥ0a�0��*k������.�t��9y�u}�����s�^��"1���G;�����f��V�z�U+�u��j��@>��Z	�_�]J/� X�|a����s��-W]Lҹ5����K���L����OT�8.#1�0yWD�f�������&7UM���iZ!\�%jl�����aM�.͆�b�dUzV]����V��d��F�-�����m퀡�[3n�2�-�4r�+iUY�1�Żi�Ў�H�����׶�M!�h�1���-���f�6�`�Eن�������b˴BhQU�Gl憥ĺ�<��Ō��K �h��n�c)��G�$�����5�S4`�Q��V1��LW�~����<��!Ц��a��؍KCR��Z\K�U+T��\�I�Æ�i{�SY��%F��| ��q�����y{ͥ	�0�DD;�k�x׾�뷞��]���UT���߾ E�z&	��)�0�6a�J��ޱwh�uT������N�W>誥~�;a��*���C�뛤{{�uk5u
U����3-wLDG��M��-4�M+��v�����ETf��*�sff8}��ԑ(� �K���0��0�r�����u�rm9�Y�w���i]�6�v���z="W-��v�wW���[�^�۵��Hnm8��4�;�_�hA�jX_�TGB��E�#9�UP�cm���"%�U.. D.�Y�EAo�Hٵ�^dn��$M�T�ӗ�K�$���}jo�\����z4����$�Cj���-bJ(ţTQ���Dz�*��u�Z�]B� �o���-���l]�;�UM+��v��a����o�b��첑� ӂ��U5�k;�YV���R���^��<�z����C͔�Pʃ:U��&c�｛�`̃����Y��W����z�8��l�BE�b3�np���8f��,t+ez�s)�}��,��f���{T���v�wUM+��~�~�P����H�����ݣ��^}V�w{.�o/P�K{z����~����Jp�	'SK9{�n�oP�CB���-�Ǽv��]<�Zނ�c��en#kyD�M�;&�s��ݽ�8�}i͐� �F+	Q��k�[���]6���ѐI�j����+�ֳ�{��sh�M������X���z�T�>����q��La�Bbb�/;�p�^���x��9�뺵���*^��}��A-u��k��Ԗl��mt��2�v�6��wZ��aڅ*C&dD!��leb;�UM+��v�v� .����.�sQ�|bI��&54/w��ַ��*��ޡU���羚�y��!CI���ӎޑ3{:k�����hgw��;X�ÑD4T@l�b��}��w�nZ;�UM+��J��{��������h��j�k*F�3&�J��w���q�'agY{�]v ���(qb6���Af��JS�'�Ac︁f	 A�����nZ9j-p�NTk��(�h�o�Ͽ�W�~�}t�؈�	JN��ݣ�<jix}����eb�^�J��u��^ G�d��"!�%)��5f+��F���uи�T���<A�ӀY�M�sy���"f={:@��}v�w�SYǡz

��0n���z�x -v��*��.n�f{�k3`E |��q
hUG��ƪ����wz�o/P�J��(6
w����SKc}T�nm
�����x�-o)	8-�(p�54����Z������v��.�L�ہ�9�K$,�)��M��]��
�v ��f���C!Z:�
��n:)<��ո�F'YwL�mN\:Cn�6%fsw�+����ZL��Z�T�Ժ
�Yh���X��ۨ^eth&��vpݝf��n������n��6֔Wj옑��Xq)t%���l�%��ɴ�3uR�mi��L�7�� 7h��3g;8ؗ63,v
ór�Z����Y��&0�5Rc��3�V��,��42]X+�������!{�լ�\�ks\W71[ڹx]ݮk�8��tt�H	<��]�e�%��;ZJ�WM`�Ec-�˪�b�������G˰G&���ͬ�P���<j����V�o�wV�����M��4�*[��/�|c;�]M#�ꩥ��+�P��}�(&
)� ���wh���SH��]׀G�R���b�מ�����M8fI�׾8���*׻�*�^mq��}�q�W��/{�!!��4ڀ�;����%J�nw`��wު�G3��x�w��$��RN! �)(! G[nJ��SX*���
��f9�t�S0�qY�+���Y��v�t�ow������%J瑽�	DB���G=�V��q�68za��J�P&gV�	6��m�BĺYcu�~�eH%d����!��#��}/��~Τ�����[�I��$#$$��r������[�bκ�sF�Ѷ����0zj�uk��*�^oX�| �}*<�>��0Ʉ�M#�޻�["W��S����h�U4��B�TB�&�M������.�f��]��5U��q��̫^�"h��LR���b�׾��z�m�z�v�
�^�wE� [,��N	C�8�Z\�m���"v�f�˥��ŁTi���0Q�lb�~�x�R9��uk5u|�}����]��S�\C�۩�w;�������b��oz�ݮ��^뷜z�A4`�Je4�����
T���]��}����2ߥR��9w��U�E@��wS-SS�fy�^
oMi]Շ�'�~۹Mj�X��}P7RD���W��d
0����g�K=ҳ:��n>��x��o�k/_ulv�7p�RzwK��`1z�W��4���Iި��2�3E�`��U'�%���x�9�׫��:�[�IN�>�ا"/��E_I16�#4#�7����k~��6�c&���]�'ttxKA�M�T�2F���/^A�F�]+\�<�q흃=�t����&=��Cvy�HB���TN��(6p��X��H���p(���;S�
�rV=��Ɲ�M�e\�ڭ��uH�FX����:$:6~�ӷ�Ї��ҥ��DJF*hn�]L��sF\K�ʾO�,Z��{Fb�\Ƈ@{�_W�>�����L��u�wgML��A�����燽��f�3��2�(�ħx-����1��,���#��U$�":�=�g ��(͸�Q�C�Ut�v�ad�&�Y�ڬ�)ⷺT�mé����xئ��7]}��l���N����� �o�6�3����e��W�����LE�;��+ѳ��̋�ꊦy�9뇼��h�I.��!��� a�F�\@o~��&#n��\m�l�g�����ˇf���3n�fj�WV�c{�"�22�Y��D��>ˆ��mY��SѸ#L�_D�D]�����ϱ��bS�,��� �&��>% �C(�I^�sr��p(�1o��&�OO�o��X3%E�E �+�B8r�E�zb�u�j��5r��^@�R	�RD� R��(�W=�n��xuo�ic �'&P	/ ��Ɇ2��v�7��t`f���*�w�j ��L/�lK�vek̈18���Z4pl��B�����eD	����-i�F�8JJLY��0��n�ˏ`������>ћ;~c0�.�a�Jѡ�����΄x��pbn�k]3����� b�N��q�g�F���̗�m�Cwx pic_K��B�/v�n�%N�������~�=�wA�ȝy�����)��CN7ӄ=���ϣR�o8��F_	YC�>/s���Dx>z޵��q�e��|�qݕ;u�)ׇ�0����ں�h����E�q�z��z���.;�t�����D[��V?T��;��tO��Y�Sר%vOm�{Yl��&��Ȅ���0�S�pZKEn�b���"p���� �Z����!��X���g����sN�~o|`�&)&��
`�f��.�ˡӾ��Ud$�I>�ŧ�Ȩ�/�9�m�Q��̖#��U�em�o��$R�R�$��s��9��ukw� e8!��Щ�| y�����5T����_�y�ŪY�LT�-l�.�^���+��*�foX��}�[���+Ȧ�����6��WG@*9���(0W8�L9��,\k�]�1���{�w��D��o{��n��L���y���2[P���oH� ���`���O�U#ٽw���zZ,��,CLR��w�]�9�U> y�fM�w�UR��Zp
Fw�>�.��뺵��B�<Q2WJm��O(��.����8���c�dt�	կ����:�۾Ι��+o����]�RF������4�~�y͝�o��3�m���d�@�6�h��\���wmsm���u�+ּ�zS	4�	'SJ�w]�{��z��=�
��ze�����L]���Ս��B͛Q����]�.1Y�t��CF+d�ӀP,4bfi�V-��
t���]�9�^ �y�޻v��Ҝ�)��i��Y�B���]���\��Y��&�N�{��B	?�v���SJ�w]�������[�B��5QAm(A�LӮ��eZ��P��woX��}�q�����s��TB�!&�Bwn�oP�����w���u�(��n��vU�!׫�)fd��B��g{_�Λo��9Q���"p��⶯�h0���z�������u�#_k��}a����X��0E�l�h���KX����@��F�F�l.6�+�*u��*�f��o��ٖ�B�ݳa�BSM��X�b��0�`+K��/YIb�:k��i���ܱ	�!fb]��D���fi���v,6����k�F巶#�]�=jƌ�"2Z�k�vw6YQs�X����[5@l�S1�}'�v%:� pt��ѭsp�PZ湭͹��;�w����1:��ޒڼ�1l�sxY����u�p�F	B�4��i1�Ɗ�v�L��0T7��图�wh�uTҽ]���'��*�oLDz"<�e�л�u���gs�.�lw�S�ݽb���f>�1����M�SK#�빵��*���z��#�L�^��YЂ`�pJe4�������t����wh�uT׾ <]�fM����JpBi�P[B��n���^ /W��G�޻�Y�)����"< ��p#��k-1�f�gFe
d��XF�4e5��(�Ԁ��,�`�-����U4�7��mv������X���ҏ�L�l���f�#��w�wXb��2�o�>����}���N���/N�w��zq����51kçlA^�o`���.�uS��?|8���xmN����VK�۔���H"ȶ�+6״k�}�l��y�� [��a�4�,4�\���L��ͱw�|1�z�m�=���ZY�:Zpl&*f���w�fZ=ު�W�w7���*�+�(s*0�	��[�4�{��g{ٕ�c�B�-��v���BPN>�r-.j�u��=`�6���U1��e3*��L��%��!4�	'sk#}T�nș�����٘�=>4�oy�B�0�e	�լ����o���wh������Ux|.���NC(a��
t���v�:xӞ�=<׮*��)*���`����طrke��wwuq 1jb���˸[�s�R�|�gg1���;&,B��-fJ1Ž`���CWUͮ\�lkr�[��\��u�h��s�D| ~���ծ��
t��p��A���O����������o��_�}�B����=����\����n)6iR7��uk���bݮ�z�ݣ��SK���y�_z M5)B�mh,5��F�Sm)��[FY�Z@قJ�neD(p�$څ�8�ޡUJ���ݮ�<|>�fNI~�]կC<<�Q4�q	�t���_��f3������URܝ5�}v�h�tDy(�m6.�{�|iR7��u��;�-�{�B�7Y�< �p\Aa��u^�ꩍ��UJ��b���}��O�#�44R��W��}�j2衋�Cb9ѥS39s*{��bq@�#]uúU�ePȊ� �އ��Z�Y����}x�{��ܿ-��������H!�Q�-���7>� �j�M:[������2Je����F�
t�>���fb;�UM,Ϊ�^�����_��a���.Xy�T݆�ؔ�X�iwcct�^щLDD8B/��1C98���X����Ɲ#}���e���W��`��'��06.����U���r�'MU+�����{�ݓ�肠�J�RBT���]գ�"_���݃.��z�ins�b
i�[J�����[����]<i׾����eZ^#���P�,8LS���b�ׇ��z�m�˕�8j�k�}^b3f�:}����(U����7�hWI�ۛ~Y��ūu���wW.�s9r�ۍ���o�ODV[�q&E��I&�
!��m�����m0�̵ՠ�V&s�гF.`�L���K��2f��:9����6��/$P����%G�S�ڌc,0��̭6]����ۨ�cu�+�sp,�d��k-�͔�r$ �	���#�����M�ec+��BbP�h[t����a�6����]4�8B��Ţ��W��V�ʋF�nnn[\ŵ��s�.���9h�K\ك��8]Sk�e3r*gkk�*�ز�e�3kVl��b�͟�7��5���z�V/>���&jI��9�U�o���R���]����^}6��,��I��i�խ��
t�;�]���3�����ީ�Y��14a��e�3����`̵���Ӥw7���>���X�Iv�}�)?�6.�^��������Y��.�x��<��-�a(A��d4���	l��F�Xqt���β���J��gL�j����h�����F�	����c�n잟UM/yDw�P��
`����l��F�".���냇���6�*�{�FGdV�<::q�W%��D�k �ꕘ�
�YJ�#آ�T�Ob�0:άz+�������\�ݮsr�wr���s�s�����{�]����H�o{��׎D(h��q���ޡU��^��-loz�Goz�����0[-4ت�}�����n���]լޡU^ ���fZ�>)È%��i����빵�����[��v�:x���d����;͈Ѥ�\��q��*b����� $v�.�҉]f�	�kV4�j2�&s̬[ޡUK���ݣ���|�N���lCAG��Jn!�6������ֺ;ާC��Ro{g�W�I�������w��3�/-�� ��b��'�Lϣ�c���iu�Վ1� 7�qe�Gy�pK�2X����Ω����j�MF�,G]^�1s\��w�KD�IA�X�k�csr��nX�9����׿~����u
��=CACn!�-&j�>�Gw��^wUR�m
���8�빥�t1�&hbwn��P���۽����t�w�o}$������0V�vh��Ё�B�њ�զk��U�c8��]n�U�U�.����oP��s6�i^���|2q�z�U%�Ї�HO�Cf��GO� M���r�dL��������%��6Sj$�ig.�۵��*�>����.ף��N�w�#�0�e
�o�|��8��0n��4��~����nG]��}ʚV�L����.�X�"�b�
������k�w<��9�CMV͹2�F�v������ko�WVv<qX�`���$m�G �?H$�	�Ke-:R�P�{�|����}{��0h��4�:�����}���h�z�i\lʞ �|�F0�Cl�m�T:`���c�.Y��X�����Y�Z��G�q\
LD&3#}��U�N�3{�������G.�>Ty�	�[f��N{�[���{6�U#��}Wx�
�ACQ�LwzD�^���}k���t7�31���0��f\>���$�guT��M{�Y���f#�yD�l�3U�<j���{��/u*�l��C"�����Ơ�K�N�Sw Iq�(O�Fqo���;#�E���(OH�n��ۭ�1%�O&�Aͽ��pp�QϷ�e�'�z��[��Ԉ����:�}Ūrpy{���2h�������]}��c��w�n�yd��;��>���t}-�`�XI��ޠ��-�I�+�-�B3�;�0�DYx3F�dG�S�h�/������x�Be��=��Nm���t\k6"�^�]7����#�Vr�Q�
�SR�TĨ�e����7�<�c�O����3*�
����_sC �9<Z]Ϡ��ܧ[�jLw\$2r�7�=8]ѡp7�a�g���摠�໰��S�\Il�T'T�$'r�t��Q������}}�
�آ:�Q������mң�q:.�/V�1��e�ݠ����s\���>�)�rbw#f��O���	\��̠�e�ۺc"ȫ�gV�ѩ��-��N�G�
�t���������Q��`��ܘ��fi>���2��-�=Oނ'tyt��ۤQ�J�[�ջ9oo��zL�ӝɅ�U�*���O9�	{����`���i�_a@};2]Z�="A޹�C��s{I�{��TF#(�ͥy���U/Fγ��Lÿ?zMa�=s��Aǰ{�騊�qn���LD_�	`^��RlB)�*�M��jKCD�f�l"�7pQ3ms�vt�!3cՖi��%�l�I
����2l#6tv,rie���T�#,n��kf��1�B5�ݛ1�j�l�i�)�k-̡�h4Ţ�Mc��6��(X�	n��������i�H(�1X��Vuu�hE�`�ZMne2:�flƽ�[6�
 E�$�6�a���V풺J%QcD�:��`K*�lz�*LE��7��i5�H�(��U�5�K-�ee���Vh�i�R{1U�Ĕ��Jv��31�����#3L�vɄ���:F�
sms36rY�����[Κ�cs�19;b��mk�t�n]�4I��٦� �*b��2رq�6%�.��$Tҥ4T���2��եA�Z�n�.]֬D��e���*35�b*鶲�Y�Fꄨŋ�V�]j���,(\c6J� em��f:	�{.�l4��%qH���%�� �f�l6�]h�F ��F��ep
8*�Ica�9���v�+�ZVbh��#�$fĳ1ik�ڭF۩�$k��V˚W����2�au$qa�u���T#v��D!�ׁ��,��݀�"�[�Z6�.�+*[�̶M�i�g0��b4ZFa��\`]��3�]�"55M,S:Ym�F�S���ЙC��%)�#L��K���c�\�&�rJ8,�s�p^5���c�. ^uV��pXh���F�j[8ˋ��Z��l.0.α4b
�a�Z�"B��0{nM�%
��1]�v�4��T�J���E����ı��#����aY���=��!0�6��h��ڸ�%j�	G9l�*�m5�jF��:*%v�+�scgE4l���]rK(Bl�2�5�j�;�������52�F�ϯ���n����97s~��N<.��W	�9p9�8���#���p��̧��S٬�5�~\���c���2�<�עn�!Ӧ5Ʌ�2ɀ�aB�0��T ��W���Y�-�f�D��c8@�}��tQ�U�2�k]���5l��.+���Zỹ[zH|w�/<��o���uJm���0R���L��ɼ6L�黸D���?!��ܠ!阮/r1������X�ۿp�_*��<��"u�سg�g���k�v���x;'e$
&m[�l˿h�N�|ݑl�)����8<��wKA�wN����l�.�n/�f|S��x8V�;r���q�Px^�6Q����ThQiZ���sc&/b(+�F"ŝCn�������:A[�'����d(�8�X:(�G{���ڡ|��5�*�ޮ|8t!���M��+=��%k�N[ymW�b���v�@�BĔx�A'��d�4��7Ñ��������+%1��H���4�E=2Q8��<_�˃+�ٸ`"��7�旺Q#C�����ld(.��A�:нJ6	�_
n��	ZX�#�7s�ө!f��jâ��5�hbg�ԱT�ri��1T��rT��s�3ΡM]5�ť�"��6��ɰ�E�m�Gj;T�.�bɮ��``Q6V
F��n�a�u)uB�tͨqv&��e�
:Q�6��\4GCZ��E�$��!H6�WB�"=��k�����:��X�i���eڤ.!ݢE|秇I����[��]�Gw��$5%O7��8X��j��@������j�9�ńp�ٳl�qYL��n�\�M#��wV�z�U,�>��}�t�GA�bd��i�խ����:}��(Tw�Ȭͪ���]�H�Y!��M
��t�����}��X�w��;�"T�Ä��(AM0�ػ�����빤s��uk7�UW��=�X��s��8�RM����4����Z�;�)���T��j��|��߹*���&���V�\E���+0A+6���A��$R�	���	��Ž�T�:�U,��>\�;��MA�!��2��[�ĸ��gҮ)D�2"wٶj�0i��[��*wRm��C��t����W�l�K�i�����H̓G;.���x��:Ns�'gw4��O�A����@"	$������i�뺵��+�v�oBa SdD]�����A�ީ��Z;�S��ϫ4ƒ�BP�@���}�9��uFoH����\ Z�޷^��H�I��i�T^oP�K�}���v�wUM#�^�މ^i6�)8�4�صYU�Wv�c.�b�4���[[���5K[\��(a6�6�{�.�tt�H�oE���^=��
t�i��yZQ��v�wUx}V�ｗV�ޡUK3z��}�c���%)BMۧC��UQy�B�c��SG�s�N����(k<6YK'z���5�B��+���pe4�.֎���1�W!k{/h����Y|(R��4X�PA����]�Cr����<~A?x��	�>�K���:�C-��M�W�v�
��ޡU�^��oz���"�-��Cb�;�D�x��i���UTnl�����c��_CpSaAA���5S2�јEL����(ؚ�ME	n�F��[M����z��ꪋ����׽�ڨ����'K	�ә���]����1���wk���x|�{�1o��i�խ��
t��u��}��w޻�G�޻�[�H�$�pY�Щ����`̵���Ӥ{7���J�>���~�
�����'<i���;XUm[�wzq�������D��w��o4�������z�}E���K-�HB[HHY�\�w;����w;��\`ZۑN�a�L
`���@��ݣ��SK��}�����
�Y��.�x}�i3��Z~0�Ay�To���]��Ir�h�u��EՎ�.ٍ��m���mC%�g#��~��Y�)�������wު�[�~,0JM��I�ͣ��+����{ݣό�Go6����!��p���	�t�����J3�����o��6���*i,΄9����P�&.��}�4��뺵���N����������P,!��������sk�}�X���ޱwh�eʋ�^�Mֈ�&�C�+���ڨR�`�E����.�v���O�E�gd����-��*�ko(�_GH��9�`����y��X72�A�ہf�c����$-j�@�����X�4s�ۉ��\��\,&��3Fa����MB֗�F�2�0���:��5vَ�n�$
�dn��Q6Ia�Gb&�W���&�v�(`�M4�;��SUF�˅���ƌ�؆�Q�і��jaIv����0���� ����д!BOF&
nwF��%�\��˜<{z�Ｐٲ8���k�g-���m��4@�.Mmi�;��c�Jd4l$���C��z=��v�X��s��|>��Ѿ�����)`�a�&LT��ޱ~ �zCM�ۺ�Ѿ�^��6���@Ǿ-��I����wު�[�w>�g��4�{�.�kO��(���U��=��ʵ��P�K�z����o�w4���2TS*'w6�oP����w��3�h��]խ�K>���sXm��-Z��H��Av�0xacrM��7Wn��e�f*!��I�&G���wh�uT�����ec>�P�����>$�Zm}wh��>�"3۲�K�FT�ܹt����rW����]��!t�_t�i�S��L�E}S�`��Og���Pkn�N�������{��r���2DGv�Η8�����s�׿�ߞ�t{�S�۽b���f7��������i��^��w��?| ���]W|e��q��e��L�n�� �w�[���*�ݪ��>|���6��A	`��i�0�4�:�U/ .�6��z�#{�׾�}�>����شRn	M�F�B�epca���yCi�	��&��0�6!�ػ��z�ilf�������wo7�*��4�(�E��-�i�;������X�KzḌY�Z o������4�\��z�U-��t7���Ofn��N�hxn-�� �M;��`Oٹ2�Z�+6��dG�2�C�^5Ԛ3�������0E���NwwN;]���F����~1�A1��O�#��]ե�r�Sd�&)׾�P��ov�idgz�o�|��n�,�$|�@�C��1wk���:^��eb��P�K6D̯ 3g�>��`�\���,	kq\ƙ�f*�4Z��Դ�� ��@�Pjn 4�ͣ�޻�G�x���޿�fx��ˍ�ȓ�P�b!�������Y=A����M#}�
���T�`��a��u4���v�:x����g��̫[��,΂���	1	�����]�#��]լު�ɞ>J,��)B��
,�Fx�m�ú���e:��9��p]*wo>��=�h�y#�kV&8���ά�3*���<��ܪ�o����JF�u�˩rsn `�\��w翿�w�ߞ?|Ϸ)E$��i�;��uk�}��bխ�2�^UM-GG��P�L/����05�W�Λe�1���R�]���6bZ\3kQM����w�.c/7��O>>�
�}���ǡ�>EC@��f1y����Csjf77޻�9�>��4��A�A�h��e6����������I��ugP�'	�Խ���{2��z\�fo]߀����N=����K�]��3g7zD�|�F޷u~�Q�����3�5�w"i�3�`�w_D����C]K��D8�m�S��ϰ�Ѫ��q�6��*9f��{0�u�cbd()�����D\vq)u����&��ء���)\jTt�����KX�+]�1Z�U�:k^��c$&�YK�%����[�&��6�1zݬ0�A�aM���ٌ�Z�u2B��"��Ưb�tҤф����SL���Pp�պ�)�B^�WYU��U6��ԙf#6�0�hܣ�.%H�m��wNtQ��s�.��i���Ҍ�:o>���F�\I���x�3�\��J4��g]�ua�Hut!��P�l0�Jp
M����񪌍�C3��}��k;�B�3��������UA����	�lo{.m�UM+ͮ7���U�`�	0�)�i�=�뺵���/}����T�;�U4�<�,�h&a����������oz�ݭ��4��|ww�*ҍ�A��n	`���K6D̯�^m����z�mު�^�i�C�\w1Pq]��cY���؏��(1K6�p�da�	��]�t����Z�]C� -�ޑ3+^i��-!:�Y�[�6)��	����(G���N[�8>��+���482�S����-'Z26oϒ�פ�������[��y�~=�߯^>��}�y��;��v�M�q��d�Ν�����çw���54�����]<k�}6߽ށL�0�-������
T�6�W����빥Ѿ����T�b`���5���`̵���Ӥww���>��X�In��>�Q�	��G;������ٓ���B������^��޷�2จ-Pp�,f6�)��R4qil�	-Ыj)�5������n���]լ���nm}�ݳ��SK܏!��A����G��W��
����wk���H�o]����O��%4P�PاK��UR7�U+�\U�4����s�`�1�;nQ�WV�F�2�v@�C��C6�tî�[�*sO��58��:�e��̛(li�gp�n���:2�:�e����ᳮ;�K&i�'��������k	?^�#G���-��5b[�''��hRZ�wJv`Rw�U�ޖ<��Ɖ�J4U},^C=Â��LZDKS�\��J��r��Vj����Æ��gvJ4�[}A����cУ �l�8��Sl�������1Ұ���"�ژ�&������L�1�r�Y��D^���&�ڼD�\���ͼ=D�qxp�+{���A�4"ţftq��o<yK'��cj�W��7��1�_N���\2f�j��7;�(L����@�k��||vd�M��t~�Էj����
�5	������:n������-bw��|�u��D��%|Vw�W���xx5�v���P���|X��sł��ux�ַ�4�6U��\N_�{ڞ���t����ۍHm@,7&���Z�����1!h�Pam�7�C��L@�E�/�V���~ɬ	��］��{b�\����mSG��� ���+޼���e�(S�=u�m(fg�5<�Q��s���͔T���{,7�B���=�ʋ`��@�U\L�vc6B��z��p�u<:�X�r�L�8TQ��Gd�
kS#>��h�b�Je�:�A��̃sp�;+�[p1ܶ�sN3����槳B{��{p��ov�{�������A�4�Ţ�&���p��p.�����T�����;eL9�w�/v4�w�!���:oq��[��5��h��f�͚Z9z�9l*�B�x@֧�* �(cF��Ƕ��,��=�]BnX��а,ٰ>?=�k�)��P=΅�>�' �	�f��x��'�w*$��sXx/��.�p|zn[n���\|��y��ۧ����ܖ��DBz?rV=�[�
����P-���X���s�y�&h����� �{d���0z\���}��\��#��p�px�k�ՕHԀu����xƥ�q-K)����[�n�����/v��qI^A���wx<o�D�w~�¹��i}�j�!NJ�o��tCp���:����Y����t`�%� #�A�B,6uѝ{I��8��%Tg�|}��E���)�!2gr�Bf��v�P	& @��Awt��ι��9%w}w���=|�w��M,g`����&m����}���xۤ{��uk#z�:�=ޱwIi�zS	8ʈP�M-��]ͯ��w�\���X����Ɲ/ ��>I�Bd��0z�ƫ\�k��a�910٪X�+\�se��
s��o2�lw�S���*�ݯ .��o�w6�����d�8b�������}���t�wz�doP�| �y����M�mCpXM�G}ꩥ���s� �}ޱsK7�b��͎�p`�0�)�J� ;�ٕh�H�*�(UT����s�x�|�������E㲦�>�s���Ol�ƺ����ߎ�%*�q��q���8�d*�l>�PY��~A8	��#����p��݈����^�|��~iC��	�i;��{z�M/ o{f/G�r�fm�Z�����i��Ɇ�i�S4�5̕Գ+��4p�1��Uı��rh�
���1n��P��ov�ilf����ec>�P����;�BF!�P�����Ƽ>�m���]Z=�ī��]��]�OtI,�a���ito�w6�oP���y��v��t�w�K��M&�n��}��
r�6�U#~ک��|�o��6���)������{�b�׀���n���]գ�"\��n;���U��uib2-v���FdK����
��gfwX��2�N��:�x����'�����p)沰�	��spl�Q@�
�D�mAA-�#m��]L7K���]����mX�+��`K6Ͳ�L��{:�[��V 0l3����l�b�1�m(]��i���w	�h��f1�D4i��fmlԤ�mB�mHA���9�34��J9M�1e:��ghU�glZE` h�3��i�⁚0�Pf�Vٵɰ���%�����v뛲�$%,�מ�5�j":+�z��AnI���X	r���<$vwj����u���΅h՞��x�����ilgu��=�C���y��UKX'�(
$D4Am�t�{���|/�P�*�Ḍ^ʭ�}V��Ƞ|MCL�[ysh��%ʫ�]��[��q�H�뺴V��Jh�BB�x�u
�F�j��F{�s~ �
r��z:4��a�л����N�����+�H�*�D̮ ÞW��W��`̻U�VV6�8��؄�`��e�J�-�p!�Cw6�7޻�G�D�U{C��woc�ƃ�oDG�l�L2�%���Uk#z����xM���H]��)K�c/]X�f�c�QX�s�nF)ܕ2R����knF	��z�+#"s.'?��柞�	��$
JH�$mIZ��d�sy�V��_��ot.c�*��	���hS��"fU�N{�����fU���
t��BG��Ya���>���sKw�wv�t�s��T�~��p`���D��4����Z��}��bݬ�2�fUM- o�8e���F�I�.�F�K���A�UG#.a%n��C\�V��L�C̬Gޑ.U\��W�>�}sl�w��ҍ�C,��%	�t�dO��U3{�SAn��wh�H�|>M�@�b0�b��G�Ɲ#{�wW��Ų�ES��R��5��CE����k\�M�B��Z9R8m\Ury�ZR�iw�ݱ�f��k�T��$i�? H �O��"#��" &�WH���m��3+dI,�a���k���q�fZ#ޑ.U\������i�Kw��%�p[jb����F�
t� �z�U#��SK3޻�^w���ϊ����],j��0��B�e�ll&B8�f͹��J7)�a&"�k6D̫��4��u�|2��w�S��}"L(dÂ�b����|[��eݣޑ.U܉��~�`悢!C ��:G{޻�Y"W�S͡S(�z�i_�x"x#��$6������z�9Y�&e\zpӣ^������W�tc�G}t��d[O^��X4�b�o-����Vm��؎�ົ��ʮ���������AX���r.����?>~��iFiQ�L48-��!K6D̯��ͻ�[����9�B����{�c�(!��0\K�cFg�m������0�ɢ9ͬe��Ԗ����(m������H��]լ��<>���^A�I��	�1~�W .�w�b��o�UR���]��M�o�#��%&m�yukyz�*Y�&}���۹���X����GE�6
M����|_o�]R���N��o]����~�j�袒>l&�p�.�gt�ǀ�{�wps�1��T���IV�1����{+#VR����Kz�r]�cw5N���2�L�I��^�����%��j�;�^eU�ȇj�u�v��C��!���I��,e���uX�5Ə�85���U��MJ1�E3�˻De�����M���B;�E�4v���"Gi��dl��۳ckX%\�W
[���Ҵ�-+cqʣ jf#�h,48�l��\#t�F�\lm��MH]m�d� �)�2U.{%Gq�@�ke�\�m�I���FU�K�-VYk�����Js���h�0�	JpZR��Kf�)uɬ.���8�Z�1�pܡ�.��^a��e�.B��e�SL�t�w��uk5u
T�d~ 
�f�j��o��p�i������^���T�=2����>�o%��)��@��*[��UH��T���o��̻G}>54���F��)������4�ͪ�W��)W}�{�wK�tI,�a���il{��mx #}^76�}B��ׇ���:O����[i}�3m�)B	ke��)�+a��9�L�UPX9�����Ѣ����~o�^�J�vЪ�ov� V�=�]ͯw�TL"S�L4�:[�B�^�s��4]�O�W���1����q�j;Nr��T�6p��X��������m�V��r��sY��9�#�g� ��$|O��lF�r�F�o~<x��
��G޺��ؽB��󷳾���80��v���SKc����|1��
q��&b�#�A	�	�1=��G�i��l�Qy�&w��ݧ1���b8d���B��{��^�z�ZZh�]T�������n]�,���4��TE�ذk��ĸ�i^�F[�[BI��PX0�0�	3j��P��ov�il{��x��|�Mo�~��bP"m�.���	��wSK�^�J�l�� �w8ֲKM����������9�%明���'�kpW#cv]٪�[
��7oF�1�G�(���$k��L��fr�1��e���x����ֽ\Lc�����ϛӅ�*1�˗5\�? � #�=ޑUH��+ב��
M�&������b�-ޡUH��T� �v�n���iC-�KHS�~�T���S�}�U4�3�)���Ͽp=�&v����lL�,M5�a0�i4�&\��Iv[�2�X:8u�g���~����ilf�:F�G�Tӿu
�^�3ɒ�,��t�����g6��Y��UH�mW}�{����pSNq	<�y�����_u
� y^6��)RĲp�e%	�u����]�9�U4�7j�y>�0��ϧUu�H�w�1s�wpq�:�Ye�1�N����Cco#7f�)��Ek�v�uf@�6��tD�tt2	$3��U�U�Qsr�;������r�������pb��F�����Ε0ov\߲D�o��0cL��t4�ca��♌�K.A(X�T�ʄ��Z8˒Ѩ�%���a���㣺T��ͩ��O���s�q�����-��`������9W��T�{���ǻ��Տ���H��S4��B��FΚ}��uS�sdK�n�z�",C��L]�����G�빴s��M{�ux���ltQLL2a�N���r�}�fЧK=�*��Z1�uIs�,��/J,z��ێE�s3.5\�^�wq�S�<�
l�i�ۃ�Gwr�C,��K�`�̣��.w!����X����4#a��7��W6���+�x˩��E{�{iZ!ѓ��U����quQ�M��eZ�T�( ����\(o�2C����3��f�͸�y &.Y<�zc�O�Iޞ(���S�v�����	q~m��I�{W�C�%�qoF'z�^X��cz�\���̜t.��g��:lWi}Fi�N]���/�qoy��W���q�BzP�K���T�dO[���:+�����۴�*�0O�,���8�\�'48=u��p]&�W>�f�4����'c,��Ѵ0]^j(e�ȼ���cFN���3�b��
�:{AS�Ij�QT�ͩfy�u�+�w=z��̜t$�ra.Q����[��2��꛱�*�,.x��.�pi�I_s��'�?���/q/�܅��
��0�TV|3��)�7�ޓ��_K��Q�6�RF!�k2�������(�S1(1��R�T��,1n��sb�w�[[q2�5k�d���:����T��kCS˫�t�����R]��%^�vR\u�)p�o����1��'�8C�N�֧X*�,;Q���Ku�F�+.,/���c��n��Vj�Ot\����	Q%�{V��4��(��9�3jf�l���~��8sU��I����T���F��'�XZ�l֪�x�ی�R���4�������8�"��e]�viJ�fˬ!�j�E�T�lQ�����Z��Єb�.#��"���w,�F$CkR��,e�1��cK,��EZ� �P�,�:�iS�L)��++b�b�=��F���c�rB�h]nSY���8��X�aa����Ʃ��˝���3���A�C(Z�����Q��]�M3����j�oTЪ�R+�5�r�˪M��kB���fl���e.��͞fIXTj�n�e�uێyk
V�a�&v����!����d���)B[����Z�sNT�8R̐�K�Rɓ��õ#e��X�DjKBe��K(�����_�ɯ���,y�%�.�%��3-!A��˂�ym�T�`6iT�cB5He*������2��Y�M�5%��͖����7�).��
�X��F]�ڈ`�Q�ct��Vm����[��׫i.[L��]Xk,х��o�C����[e��[�Q1�@К�[*�3Є��X�Dv�\8 �R�:nF9�ۀ�"WM3X�f�.�1
�X��;Sp�-�arB(כ 3meM��v�üw�'�0�����W�t�f+��%�е�a�+�K�%J�b��b�ǰ��h���.��%��
e���$Z�[m�
�e�Vj�7�<M�&��j=\=���kn�� �0��:�f�a���f��]�U�^k,3�,��8c6�1Gf��3W0i�sP��r��4ʴ���g]�i������Yj�,Kf; Ħ�1��B�iS��$Д��4��	%mW33��8Vh���L�1mHM7hn%%
	v������F`�Y�&+pMK�L��LF��l2+l	�i��܌�`5V�]MHIKP�(3�,~t�~}�������h��N��v�K�"uM����ä�*���O 716h!|mCq��&�O����K��n��(�enG�mA�k�qs��jf@��ΚGM�j�K4��p!� ����3���������@S9��һnd��H�R����L����y��!�ݢD+ F��pd+V<B�)�b�r�'�����Tu׋ ��JI^w�g-P�f�3��m������$�5w��PEiV\�j�z-�sV�Nx-�+�1T��T캖=TM1��bޓ3������=���������zFi��$��
ʜ"�eVQ��
3�a�t��=�{ϝ�|e�}��x�Cܝ�;�ώQI������@���DtI�[G)�grJ�n�����[�LZ�$$K�0^�W�6�7K:C��>�9�yъ���&��2g���GŎ��rf�o�r�{o�<C�g�G�`k�RǑ��A#s{HӀ=}����c�w�ZviN�u��Eۆ5�b5�[�x�y�l>+60�-�׎���t���D�@�qbcIx��w~�gsG���Q��[z��7j`ǂ)��!RV�E�6@-����h��M����J@���* ��V�A��ͫy�,qx�r�t��0�Y�_!��`n�*�jB7KQ �^6���cv-k�e��]Wb��ֳl�bi�0�X� ��Ke���k��s�᫐��G%�\�rʱ�E�ҳ^u4��̆�`٥:�m�����b�K\�ԉ;��,)�&��;�wQ�1y�t��w	�Kw�f�rR͙u�º`WZm���3C0K��݊�����C��C/�M���
�W�\n�lt����\�9�)Fƈ�L4!�Y��C�����.��멥��z�m�^�V�O}� b(8�ػ����IE����͡NV{hUR�s���&����|�{�̛G}�4�6��߀y�ٷK��<��8 �`��h�H�+��v�ݣ�ꩥ������G��5�4�3���fu���6�n
��1�	�����ict�u�#v�V2�ˢ�9g矛����ݭ��4�ί�}�ճ�"\��ڃ��'��v�{��=��_�����8MlUɚ���vpiސ����4�9�F���YEƞ=41NИI�*n�)��t��>��"� � �$}���,]�Tqݺgv�ʸE���-�4�}����篞�B������}��<iy�Bm2Ji�t�益�͑/�g�]R9Y�0�jP�8�	�����\���X����Ɲ{���]�%��q	��e�	�t�=B��� Fw]ͮ�w�����4�����״��v`R�#IJᦲ!�4s�2�v�7b�*�-6�#ZP���B0�i��]�t�gUM+��}sow�*�-ց�SQ6�4�M-�o]�}�c�z�U,����[<k������%��Ka�@m�ͭ��
t���T0�Du���cݘ��KHu��'c62��.[�]��������8���
b�n�&vy�;}I�f9]��X7z�l�{�{mMk:=�[��0"22��劢ƃr��X�)Ђ~�� |H'����ѝ�sk��6R)8,�LTׇ����fZ���Ӥw;�������X�K�y�DX�����s��ix|.��'��*�^oX���M>�}�Lئ��1nRjbh[�R�X7dx,بi��l��c\��J��B��������wV�7�S���<>v�wUM-��
<�1��-���{z�{y��v��t��u߾�=�|�Mh��6)���T���O| �w�w4�oP���G��a��b����z�m�=���Z�ޡN����4=���bq����)�GB�x�F�Tc�l.ȸw��thJ�������<w\���:!��7uGo���=N�����_%���An��N� �:Ka,���>XEYlm�[�����\ܷ#����^��-g�`KBa�I��G;j����;z�ͬ����]<i��{}!/�p��`E��a4�ZiQ�Ԩ6RQn#��l-�m��ZF�fO2�lw�S���*�ݯ ճ�ꩥ�T��M�[d�ة�y��~}���t�oz�d��>�y��(D����6h]�;�UM#��S�>�{z��,����Yf8�!6�$�Lү|>q��̫[��n�
����w4���6��N0�����4�>��`���)�H�o]ե�wc�k�YR-�h���Vrf�N��n�Onj��y��r�;t�3Z�u�HJ毮9m,�Blؕ*��nU�'T��y���b����:�G_"�&-ܮfɋ)��5�6�|���,�u�8.a��+6VhK������J`��ۛvQ!nWHQ1�X�x�q{F�T���V)K�љ�\Ԯ�Vn#M-���Y�2���it%S0h�s�
�7`i���)[�1r$غ�c�X��.4Lm5�La6���V���Bȍ���5t&~�ƪ+yWKp�����1��n�G97$�]	`ú��6�xp��,�#4&�	(�^Ԏ��6�.%`�E���G�in!����*�/��T���M#�6�}��V�oP���x��!a���b��r�4�����eխ��
b��С��և��pN���o:�GshT� [��`˵�)�K�x�66��wW� z��-���T���Mp�{��o:a��pKd��M+����^��:�h�����F�
t���<���BiA�aB��m�z���]c[�X�JqW�W_ͮϐ���G6*���K�67u���i�Gsh~�}uo7�URֵ8AM80�f!�J��o]�μ�{�qs.�|n�B}A�b�vs�r�-;H�z�r��=!nt�;�k��jf�ޓ�g�L&1UǤ�p�\�jq~b;�ݵ�8�8�#*�$�����.�e�]ݹ\ � �A$DT]ЧJ��*�ݪ�>o<�B�(E�d��.�w�TҼ�^�}ʸڤw�뺵�C�AMh��6)׀�����G;�������q��.i/w80���8B��w)�J���w�+�z�:[�B���b��`��dõ�G9�f��h��[X��T�F�cv��2��&a��h$�ͬٙ�r�M+���>��ܧ�*^�:=�F6��Z�ޡ^�+��L���so~Lݘ��#	Ce�ZlL��dL�bx`_<��m�"�L>�˺�2�#�ő�5�c1X;�����ͫ�{����w����Fؾ��Ҝ��3��b.�\�wQ���w7w]�`�`$	�SU��ޡU�d�����m
�}�
3ާ>͙�@��
��>~ޱwK!��Bn�a�iR;�뺵�>�~�j�oP��ov�it�}{�߹`��)m��6ŭ!krl�e&؍�4\�Ll��E�H��m�!����+�z�M-͡UH����4��z�-�^" $S��I�T�6�{���9�u4�ffQ���|[|{���	��.�|e�9��u���/X�K��URV�&[PӀ�u5� o]�#��*i{6�U;��׀�ЮН�Yp�f߮�mt2y�f��0�3���G!p�EFUͣbf]��7W�ΐvz�l�����PJW+~�6u�t�w\)!r8�t�v⦋�莮rtŤ:� ~��������w�MGF��f��J���n���G;����z��x}&���}�s�� �YG#-3�#ge�ю�V�sJ�4ڊ����X��ߞ��ߟ}�wh��.Q�Ϳ|>�[��Q�z<��6*��t��|>���U���T^�P� ]���P>�6�!0�7N���]լ��){ﾷ��.�W�9�AH��%�6���>=ޱsK;�b��צ\�|���ʵ�x�(h(`��b�,͡UK�}�w6�{�wV�oP������N�&wv�_����W���lM
�_�Ceē��N��Ƚ�K���'E\�'�����uwFu�]M�i]W�&�6��̈́�a�n\���JCL=vv���u&U�ɥl�����	�I{�]�JF0ԫ5�4�rs�ƽ�eH��\�U����[HgM����珌�G֘�aK/a�"��2ۛu�J��ŵ�MA@���f��[��Ֆ)���U�I��DعM+�m���H�Q�:�#��sH\G�5���q���:���� �B����P%��)-)�a,),����5�ђ9��4��bM��,%f�Ժ��1��CVjJͭ����D&�B,8lO�Gό�G36�do���\���T�d�"L	a��(�M#�޻��x���T���]ݎZ_��J��F�XpἻ���1w�U��ު���z�㴦8$`$�H�m��������sfs3f��f��M�����PmU�n}�����;�P��y�b�֞�H�[�߹�&�m�l4)i��M+�+6�r��+"�h���Sd�v5��M���ׯ=?�B�+���*��ݪ�[�Z��~-�I;��s��xs�"�"�}�j�.V��)R�r򚽃����WǴ�r��ZG�	��R�/���M�y���w{|���g$W�W��7߻i��c��.t읺v��ܺ�r�r�W]�I����S����?�_/�>xk�(��W��U��|�

p�(LS���*�ݪ��l��ٗ|�q����D&�m@i;��>����Ϊ���HS� �w��%�P��eÇI����u������P����Qq��u�������n�i��Gv�hM��E)��Kl�U�e.3�L�AA��8l��3{�*�3deR7�^�}uo�}빵��P�L@l�LTҽޱ~ ����H���i\fЮ鷓��$T\�wc}降�����GpB�h�˩hVD	g=�l�o���m�W42MK��b��2�wi**P-��uإV���c{"΍0vS�2m,*����Q�/�Y8)n�ws�Wq��ģʑ��i\�^rqm%wٗj��%ǮT躼�UuHUƪ�Yr��u�"��kQy���P1��c�+�ºH:'nnUl�S�w�0�l9�D���ͼ��[K�]�	옋�c6�C��$�9��oh';�֓q��.�cP[Q$�n XJ6G�b+6&���_��Y����M	۲�I_�[�����{�9�q�U��~��)=0��{���I�
g�b:��x���U>�m�y�:�����	5�(7�1��H�W:/*+v]H'y-�B�<���tO�[g�*�|�8�w�(`���_f�Q;����u����d��r`�nм0{��拣6�o���;��ϼm+&9r����p.E�D#�o6"&�\֛g%�NhXv�D��W�����+�jv~5���-#�!�ހڳ�:��%(��k ŗ����+N[�?*�=�{^.��:����nr�n��޼n%lD2cMA�z�%��S�R��u��A�][��uN��J�^`��P���}����l�$��n'�I�]�ov�w����A��(^�.ozx�j�i�
�N�uEU�a�/1ur/n&+pupq�ES0�9Hn:��8�پ�Y����|=�K�����x�8,�{L�4�Lng�F��׺�<��M�1�{�T|�nt���>���S��䳐ُGI�{d}o��
���1�`�5N�E������ʴ���\+��^������ 94�.�.�n�H�/��$���	���8V�4NL X�в��Z�Yd�����L��G��SY,	aW�u|�.�G� בf��-�*���D�(���T/ex X�Q=��/&0`�<��O"->���W�$���d�Ԥ-�V�������F�:��P�\Pێ�kp��b�H���x��8@_�ē����4��vUO��͜7~��ռOLj�}ۖ�͇i�;��	��UD����8껕���pV�X1"Av�?��I�q�'7J�n�����vwE�H�d�˛5j�U�E�����»ۭ��4j�`��,4\��ܣ{b<���G)��R^9<�I�ѧ��#�C#w���_F��5�fmdab��b,�f$�P��;x�^�����r��wN�m��}�_l?{�x���ʃg���ݞ�5#�؍ܾ�r����/��Y-�.d�sN�	�.�3���E��Ȑ 0I'�;�A�f�u��E�&%��CfW��_{�NF�)�͙���uT�{xG��R1%�m�ͣ��*i{��o{f.�T���M/��N�i�V��2�HK��&nb��l�e�8v�hXT�u��҄ڂ�M�l[���*�ݪ�[޿|V3��
�K��E��ػ����x}�}Y�)ҽڮ ��1ȓ�`�����w��wK����z�qg/#DAB/♃
�p ,^���wH���ڪ��ǔiuQ!�{�х�2��T�&�]�B�5�P5���*��Z����Np1[�M^�wp��9�����T��R$�t�/ �1D�f�v�c�]ݺnWt]���˻�v\\�nN����R@�%:���������|�2Э��W��*�x 9OT�gUM+�m
t��I��,���DI���h��,	M�����q�u�;��&P�AB&0�D0�����SK{z�ͣ��<>V�{�.�l8�/4!&��*���^��dwPS��T/vg����AM�Q]��zC����w���=JFv�UD^�(�b�
^�|���L�9�ڪ����X���G�ф�6�CLUFGl��� s���7ޑ3�"f==ұ��*Xd߼��i����Ρ�s-"g&B�A���w����!��v�3mp��î�Ot�5S�qT�l><J;���뫽!��
"P�i�0��"2�f-��tjfhe��X�` �u�\���I��&s�`�K+3��eGMb�t�պ�)c*R�5����d�:�+	�@���y��1O-��bbmj��X�+Y�sN!L�3V
f�\�h�K�ln�j�4k�5YCf�+)pdl;Q�mG��5h��k����{��%ۛ�5˗M�6B�\�s]9�%�9��Yo�;����&K,`��e-�R�u[SSk�8�բ:��<���]�L����׿~�TvwP������{1�>2�v���1	�����G�"|>i�튪G=�SKٵ^���w1p�BM���1SK7�b����+�L�wfU��H�*��-i$J.
�ػ� 8�z�i{z��ݡS]��<���^k�({��L��%�J��^���
t�v�U#~ک��}��tyy�Dz��anh�:̤2�����֦hf�ڎ�cA*A4%����B������[O��SU��wq��"�8��p�D�^uC����^�7uKo����޺�4O����MU_o��ε�uRr�H�Lt������w)�W=�W���ߟr�����p���-��vup�أÜ�;�+��쪙��L�̑��K�{Ń��$��w|W��ۺ���zD���U/<y�`&��%�u5�|�����4�7�.��|����%�
&����Z<�Mx|.��ݣ�ꩥ�ڪ����>�_�Tm��jT&�j��n�[��[P�n�2�v��¸�L6\4[,$`�-6.mf��]��Sƕ#��~�g�4�^P)A�h�SB����W� Z�uL��ީ���
��[�����LҤw{�uk#�J�4<�'m,X��v�7��8>����4Ș��Fp�;��]��D�R:�HI�T��6��i����YQ1Q�����w]ݮ��wvb6( ~ A�<z�j�nt���6;⛆�'w~�Ps��]�t>2���+��f\F�ǘE�a4�$�LfgUW��ު����wp{zC����1އ�_4�BU�,+��)C]e�.��͕��eZ�W�[�s��a6�4�f/yO�*Gsz�doP��}so��URQ�������i:�[޻��V3����Y��v���|>v��`z~(8)���˫[��)R��^�}l�u����z�mws��)6�2��Mx|w{e��5�J��޻��n����(�?tE�ݗ�{���c^�ʤloF[+m����)�Q��v$�@BK��g��������k�&")(9n� {�˖~0~@wr�ỻr�K&@���3�)R�
0\�wh�uTǾv{���}�'w�U���!0B˛ش���s.��9a�4ef0�l�a��f�i�P�L��l�٥��]�f��ʖ������ꩥ��|T�S�a�w6�l���	�{�*�ll�Ӥs��~��F<c�6���jb�.ޡUH��T��[��{2mt�r��kpb8p
a�]�}��W��G��SJ�m
U�}���t��k�j &�����u������P�K3hUR���K��\����S~�<gs�kN������͚o�:(��QU�;���*բoJw��ݼ(����{��I��о�Ơ���[��6�WUr�&H-���k�����M���ۡ�#�ٰ�[Y��e��b�%&���U�-m�Z�\�RY��V鳶T.��~>y�1/��&�f�L��J�e�*���h��D\Y�S�p�j#
9���T�3K�-b2�����5ځ�J3�ia�葮&62\573iwQS�I�����s\Rg:wt9^��/�&=_K�u�ǮWlf�*��^u@̦�6�h:l�+ë,t�UA�������)R��T��������޻���d?"E�HS���+�}�����N������m
�ow�(D���,��ݍ��f6�z��}�#e��VzjM���Q)3+� /oUu,���nm
��q��sKw�@����4�'wV�l�r���nm���ܧƕ+ͪ�^ ���6�#��ۚE7\���Bh�/4�m���j癦�]b�-��8L[���*�ݪ�G}�~���t�r��rn$Xi���ݭ�>4���]\}A����U}]������θ��uCzf��j�UU���]�'��&�%�wP�[�s+�#"> � �@��Ę�	���`����{�K���+� .�5��G"�mÀ�s4�����=�%� )�m�˵��eJ���:
�H$��� w�S���*���Mw�>������pi��M��-1SKsk�ݯ| �<iR7�U4�zD�]���}�D@�h���7�nl&0m0Dٕ[�ME��-���Pλ7@A(pX,8c3��3��Usdx�����w�8%�&Kd�\̨���}��zBq��UH߶�� U��@P
LBYsh��B��f���:�*���{,O��q1�WTl�p)�)��r3跓2v���7�|iMтuWXi���z?=_~�� xB�-���'���򕑞۹��wB�[.a�4)׀�>ޱwH�uT��ڪ� �b�?w�'l�a�wka�+��gvd���R��U.��o��bJ%�kMl���Ԋ��Ī\���n��v���	EÆ,6�i�8n��wUU#��*i{6��}�f?yO�*[����_ͷ;��w�O��M=ͱUC=�3�3� )fB
h��b�����C�+�|�w�̸���j��@:a8)������U1��=H�m
��?���ͨW��.Tl��昘�\"'���abͦ��3�F���f��2'd�P`�i�dNZ��~��%����=�f1��� �^,�(B�����>|�������c�|وP�D��*[�w6���;�)���T��j����xO�	�	$�C������\�v�`�����f���S6Mɳ3n���G}�4���]��S���-���z�m-����4��R�����^F�hW [��y�(,4ۀ�b��yO�*Gsz����U9GwhT�Q��Q`�ڀ�:��~9�!�Vg�w~���|iG�� |
�H6��Z;�%�~ n��G�2�{2��T3��� �H�$ �m��ַ]_ڶȨ��?h��hu�����x���l�{��g����fL �h�$�*$��"�U����5���U͵[P�袨Z �""o;����b��Z��j��Jڨ!YB@QP�q.��   f*���kQ�� �y"�Ƞ����"�� $��x
"�� � �"�b-�����b���
� f
h����e?��v>�\̀�h��?lTD�TTP���6>7�����{�_S������������������)���O�?'��p���+���8���S�?����=���~��?���j�e���~�'�&��@U����!�^O�����t?� U�*#��X�>�1�����|?�����K����_���O�!������U�D�����"|�m?�G�@�3��)k�h��!b��7�0�Kg:�u[�?$��P�L~o~7� �:���B*Q��fښ�jm6ԳmKEB,T"�B+`1��V+`��B
�B�P�T AX��UZm�m6ԭ*��ښm�fڛ6Բ�&ږm�DT 1P�P��B�B"@
EB E
AX�`�@"!(D#)���$T��jT�R�mJm��mA"���`	�$�DVԶkR�kM���)jeR�ښ�mR������D��H(0D��H �D�#H��#H�"D�Q"#H"E �D�H��(�֕�6��ԵKV�ZR�  ��"�F*�Q"D� E !H*Q "_���EB(� H�E@b�A�$F(�(�A�@ ���X�DD�$Q"� H�A(�B
B(�����mJ��6�ͳkD�Db��$��P�i��ҩmM����U�����Z��kKY��SkAH�D�A(�P�$@`�H��A �0Q"�*P"!H�EB(@�T � ��EX�DH�@���mR�YiMR��VSm)���KZR�SU� `)�EB�U�$T�EP���E �$H�E�$ X�AP"��$E@X�D+ U�TP�$A@�$AV�U�A b�F(�U"�"E(�@�$�$D�$A�$�$P�$�$(��F�m5�Zj�jU+i���S[6�j[-��kKT�D�$U"�b��AX�@B(�T��T"�H�D(�T�$P`��A@�$�E�$H�@�TH�@�$A(� "@ )(��$@�E�V(�im�SV�SkMe�+$HQ �D�H1D�D4Ҷ��қZZmi���*�R�56�ʩ��T�,����YJSe4���-))(���)��QL������Q��&�b�*6�K"������΁k-�������~��=O��]�qTTG�C*0a�?/�>a��a�����'���ͣ�x6�>�#�:������|HlU����ҿ?���>����:O�~%���Ї�7��G/�.�\�Џ��N��o������U���? �w�����?G9����������~�@�?�U���֌_�e�y�����C��������y�8|� 
�9���F+�"�#��.�����@�>W{v̰�Զ@2���7������*#/�?�~?��P�_��*���u��A�C�h����~�����f3�c���e��>/����c�� '�X������]U��C���o�ED~c��#�=6wc����p�$a�`�?�d/k��fq���[������>���>*n�n�ߏ�g�`��N�b���O�|ߟ�kC��>,�^����~�8U��d ���ϛa�3��~ܨ|���`��#�a�@}�!���������TTG�|�%�n�_����|��˄��}]�A����s��/�3���y�Ȼ�)��qb�