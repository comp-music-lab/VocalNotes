BZh91AY&SYʒ*�,_�py����������`����           �  J�PHRTQA*�A o�����  R� � 
�w�>�V��N<�M6��y1B��Ӷ�yc�P�D �P�|s�r4m��sig��ow�<� �jݍ�
>�	wQS����������k�sǞ�ӭ�:ww�T3
QG�$�e#���ٯT�B���=+َ�}/�A!V:)�=��e�hU�Ǐ=ގ�Yc��Ϟ�ϸ�E$��4;�IJ=hև1�t�h�z� :���:q^�*��x��P�l��+�I@�r8�u��\��iTH<J�tU ��9�(R�֎1���P�b��"RAI��b�;�U+M��.�u =i� @     S��)A��1���� ����R M�  &FCLO�*�JzmH��     5?"�2U*0L  ���d� OI�T�O�#&&�� � M4`���	�U4=4�S�'�1��2z���0j���>�i�
�QAB�^�D8��� (X���� ��X��*��@#Q?�}�R��p���5��J`���E�O�>�����Ј��X���:�}���E����Qn���c|-���:��\����^%�Y��ݰp_ml�xl���m�5�-E�h���xh����h͵]1Wa,���7qs�������Ȑ�٪�����F�Û�I0�3e�^�\�јxc�v̩M�t��U����;�k���n;�8���j��a%�y���s3a�������X�y6�hj� rG�QWnӛ�'9�P)�Sb`<&ږ��r&7����>T��)����ә:�qc�(r��`aiDs�uM<�Un����M�mr��+�z�gK+K�Ul�z�k{`�T�^̩wS�;����M>Gd7�q��qi���J���3���a΄�KM��q�iR���=&*o��8�����'-�7r��hvwq#�Y���;qw ��`n�br��p瓶�^0,���su�xC�^�坿Υ���b8��U��Tl%:�ވ0d�ĮK��Y�.7]����m�ᇧZ"�tb����K@�1ogV�Gp���I[L6Տpp5��g�K%{�jT8qlb9.Bn=ulM��H�}�
�
����E+-w`���b���#�w�����r�ݭG�i�s����;�a7�ޑX͝ٸ�ѷ�q�����|�, �<����x�bq�YH]�ZUcx���Λ@�U�D��^'��ݣ�����[4��y�M�-KHU���}��AVL�Ҧ�mly.��v\9�7���)^��B�U�@�iIX]TP�Ih$��]�zkbgQ2q����-,��!N׃Q0�,�p����p�r絝��X&�:��*��2s�.��7�ѣ,5��T�K�����{Jܸ�s�)�i����̀/n�.�	IG����83�<J=eg�m~�|(�la���Ӯ�Ms��\�8M�͋��]c����{��x�q��噽A:��X���O#�I��<ݣ.)65���IFL����˲,X��0̚qM8%%�Nw�)a�����#��G
g0n}�WET�C<�.m h�zb�W$��g �;�.��6K�2`T�����t�*�l�LV��M�	�F�s_-���'�7W��0ս0�ys��+�-[U�y�(�wm��FQ��N�929��q�EY��<���::�[$dE-߯of�v�׈�և���yJNr��.�/j�'w��ԯ6ZՆ�٨��.��7�ƺ`�n�������ԷGk�eW#�{5"s^��ݛ�7#l��f����Z>Ѱ�aB���h� ��Cin�%=i�dt�x��(v��a�Y�.�߬E��{\g���s���96{&�s5��4��͜�47�hۮW�WMߧg>����sNs�����
�6|����%�����	n7�Gc�^k�W1�u���3��7S�G�r-�������,���{c,�����{n�@�rp�ʜi��E
�����zQm��q5�qCO^�Ѷ���i��Ϯ ~�H�&�8p��p�\�5���vnT�N)1����/l�ҬC\�h�Բ��I���*Xa>�yǮ��F=�hTF�#���]*�21�PVlѝ�殍�=:r���'�B�Ӆ��t,���q��8���W��zB���Rsn涕�f(g(�}����˸ݔ�.tkN��F���b�OqyV���Op$� ��g(�p[۰���PE�#�`���D'x@����+���Q�4s'2UǞJ�n�F�v|쁻�3��!�-���ʫjig%��J���	��oIݦ��f�`�3���C�����Z*I�q*��"�xB�gz�;w)�*ud?��jHr�[�9�� ��8LT3�vv��7�!"��3�:���G0�)�X�:�'+�A-ee�)�J���s��DX>x��N�W*5���HF`�ȸf��7f��I��K!Qb����q$C�gbu�Ȫ6e�]\5��4^�^�2v����G]%�4��Z���t-I��m�4H܂lKn<���*����p�w{��˪\��{�T5͂�C;Y���;a�	��O��:��$�Ԏ)O�M,d;:�lS9�����ɝ��J�l���#7���b=��ӊױ8v�d�7�v�j9ܤ���]������_7��}��1�ðL;�m��bx\����=/����H^Sw�FшR,�>>�Vӭmnx��m;�O��suY���>_y���{��?ӯW�c����^��Q��!Q�>�ۿq��a��=�����^0gK�4�:��W�l69��Q�����θ&�'�!6*�6�뮸�#u�ZN�2׬����#��e�˧��y)�����$�>��7jG��k�6��Hۜ� ��r<\�a�.�(�s����|㮨�M��#�婃���M���g�%�6��<޴��\����|�7]'mk�h[��B�u��\����Z2��\q�vkƎ۶�(�8����"|��"+��D�뛮���.ѕࡪ��s�=����ũ]������#s"6}�ݻm�L�	ZM����7���g����']��㷥������\ѵE��'-�*�a�eּ,vj���t���W�la�j��t�2]f�{F�k�=����9����P�H
&��ڃ���TŞ��]h�a
h�.�k�KU�poqΠkeoN���i�xr,Ŏ��ci%NW�W�E�m��a�	��f��0�0�606Rh>uzӨ��[�^3�u��ڇ��O=��]�K�����fL'#��\Jn�6h0B��/OW��6�Rq1���`��b�v.�;����Bh���:牫�ٲ���Mu����{E[ѫv9����B�a�� ''^�hY=�;����:Ц�)�!,�1�#.���]���/E��m�"�S��@m����e"��eVs�C�ǵm\L�Pi��7��'��/[�j��g���x)��ͷU�:;�y\u��3��Ll�7Ew\˦0�改Į]�Χ۬糺��O���4�<�Ѵ��Q7���1�nX�B��4����]�kf�}Y�M��[m�ـ$Ԍu��6^�ۀH��o�`>|�����؍"� �]ӄ�b? y�۪�:|%�T�e^�1'T�n���v�]��^�uS�u���g����RuSP�՝)�\�QKt͎f#�D��1q��ΖC�6���6n�ڷg�ND���s�d:ܑb�u\g/ )pa�A�uX�Z�!�"R�Z�9yG�r�-ت��U��v��y�Hv���^��eH�9y棲{m����8'|b{]���智yp����v�W�G>����zyp���K��K1(�#��B2�36���Va��:0v�qѽ��S�ٖ;8�fP�E��D���f:��gr�Uj�����	Di8�فS����2�ɧ�m�:-vw9m	����sOF��=��vb��a�Nx�j٠n�,Sr�g��q���b8��m/3��F�/W:�sx�s#��Fl���f�d�l�CYl׷��zֲưBMt{�s�g�۴g=�g�X�0|ώ*ѹ�*�. n��S�Z�k�r�+xu a&lN�� 
[	����'K�7W<�[�
�Ӫɋ�V�%�,r��UxD��ƪ�"k��dܡ���G����δ��cV-p$8l���M#�ݱ���sȩ����#Q+�u�һ���1	����P�e	�۷ ۑ���8�WRs��+3]�M@q]�R�Wh�Wn72Ǘ���M0bqs�������ʝ��k�}�Y�2���|Ż4������Z�$tj�g��u�:��p{U�u�mi�)$`��t���6C��<J�7GX�e�܅�EmΙ�]V��wܽ�&_�P@P�| b�A	�u[Ȕ��Ux����K��~!�����Wg�$��_/s��n吹_T=�cW��۶]���Q�2�*Y����{p{�y�B�DѰE����<�D����Ԃ8, z���{��G���N�>�ޑ�NV�W�BU��v�^8�pZ��2�^�d�z�30!�*�k��S�XK�SZ;�{�fU����Á��q�!J����1���=�%����Z�v�n����X�IܿJ8T�F�FV��ףMl]�pM�ه9d�÷o.u`�{��.��cܲ1��3GvzX�e��6w�{�œ�Ak���h�]v���͝�E��`��Om�h!�z%�� wͦ��tz6�wO^�w�ݏ�]�n��8����,W�����v����}��H\.���eb�6{N�f���zŲ�!uB2���u[��uy�M��𻝜�:Î.]��t���IN���k}�W��vC���m����HB�d��c<|��s�M[}|��d�C��n�N�Ǻ���}���M��o+[��,��Z�ٚ,��;ȆHW�f�X
�
����z0�7��h���JB��@��=�"�E<=� X��d:�h>#C=�w��M�}V�2cO���h/�^O �]���W��\SK&,wd�XD�H5��h���6&H��>�0/@wg[��~����"���sv{���cy��n)�S�)V��N������4�Z}�G{�v�W�s �c�]�u��9Q�2������yٚv��	��#5i�ܺ���W�,�](gތs���gd�W�Fvs�g���J�^��n���C����shN�6V�%������!P���"�8@G%�t>��b����OM+/��'�ǌ{$ync�/��!��OH2ud�;��G��S�t��m\�9��.y	A����ѧ�/�d��8�J�r��벷^ҳ��W�̷[Kv��z���>J�Gy�,�݋G`�g��za;;43p�$�՝xKC|S����� ��u+ٯ,�IPSx��Y��|�S<=o��-i�ߨ�w�7����qf��{(��X���b�n�l�V�H���g'���%e���4���:(�S���7K��sXA�!%��rd��wF��<}5��F-MF���]��,ST�O��"���>�|�ǅ֕�TX�w&�%M�
���՞���� =�쨞��Mq�r�2�ޱŞ�:�m��� ;�Y>`�N��T���)vD_Q����=� A�����׀�%�^�\7�D��zC�v��л}�sڱ�Eȩ�p\1��m�p- ��p?��}=�w�jeD�q�u2CzSܭ�V��DĤF���\tyG�=��CJ>�3˺G�I������	�zN엎�XgR���x!>xn���W�����|�W�c�3r�+��������w����0�=�����O��5b;��t�4b�w�)�W=�_;1���,3��@i-�m�x�c�1��@Vh��VG��T�V;��s���Z6�rg>{��s���{�`o�K7t�x1�sݾ���N��7_�l��%�O�u����=����C��k׽�j��O���Gu.U�sW�~���8,s�R����T�\�B�F�=��n_R�U�7�/k���l��;�f�A�o��A���[E@k4��q�	�r�<�w�v���{��<o�w.�H�;ݳ�z� �MX�m���/tN[�]ɝ�=4H��w�e$&���[[�*idp��W˸U��tt�Lm/{���uӻ������M�-_���#�AE4�I�w婍y�F���O��i⟱�lP[n��0��T��k/ ;���n�k@x]���/{�����p�����W�Ű�ُ �m;�h��{5={��I݃|�<�
����x���G�p�!��n{|��˪�e�h��Y�j�ٷ <�^����`��^�ANΜiDhv2nACpQ`�szi�!I�;4�KP�x�ٽ��^�����F{X~�'
N�����u�'�iy�.�|�+;�ځQ���gܔն�E���s���='������� G%���������5�!q��^.Ĺ��';��{����=���@>�=��s���L�[\w�z�f�ɜw�1ȹ���3��l�[Q��ō����x�?����O��L��s�iL�Ђ������P�AF=�ºP�:��{�R�󦮞��8������(@�	_�&�/��^�}$}ϙ�|�21e�f]�*�󫘗�p�)Ɲ\�V��GF�	s׋��8��Krv�im�)�[�<>�S���75�nkui�̏����N{���^Q �������$^�\��q��,Y��y�x�
Pxu�Y�JB�n�ܶ0�ݎ(N.�^��z=O�Y���:��6n�Y�ZM3l+4p�\@H	��n4z98Ƽ��G-۞��q�`��r�6��i��+G.s&5�u+���lʌ��8��[�`�nW�4q�m
ǗV͸G�6���"�u�	�F�I��ÓA��Z�\�Y�ux�_7Y�-�>���E�y�cR�7nG2�?���V���ھa�a�$=��%-W�o|V�
��дC�w>N�������r��hVpJ���Fs�ŵț�90u�gE��̩f�b��D�y�k#e�t��{�h�z
��ܫwό�y�\�ˉ��T��D*W��#^�ٜ���d��r�vsq*�@T;�;�+*�W��,���|���4�ڮL�&Y����|�z��C�u[�qgQ|�Q}���_|_|�!���CT�%�1����d�]`�9���[r+�<]�dH��vak���ֹ��4gr|̴ecʬ������s�����e�F2Ķ��P�����Ǽ��񠂍7��l�>���C��d�"�H�M����5�I�|	=����S�ܞ��~	��8�h��B2�a(vR�u�-��[��#�S�rv{j�pRܽ�%�!E���a�D��	)k,L�<�7�v�S�¿w1��)*�ʱ�� 4_����!����^� ���D�2}��*0��I���B�q�fz�}�.  �[E�������ٖ$��ܷFeoO%V���p[*	q�
�*�1�K��u8�,���ӟV��*�#)�W�����m����.P�#���G��>?y>ux�i��ž�"�q�np!A)C*
!WTwh�ͨ��АX=y�����B��:p҅4�F<�r�2lK���`bF.��N���N�P��B�h�E6<��$4
^�>!"�!��:�X*r��Ђ/�g�L655Ќ\��)�ȇ�^�g�g���Q����C�꜎E4��L��!�m򜈈S~<n�r��촮<p;�ꪛ���gcPs*���2P�='u��'M�ӷ��
�h��׊q�bY��lҐ�Rf��GiBh㍞̻t��)Ѯ� ࢕=s��l���k�ь\���[N �� r�V�%���Α��x^8���E�fq�̱R�ya�R2F�x1'ef* ��7�͙7�"�P��q͡ҫ�+�]���{�Q��:�Z���6�%pԮ�f�.4k�ׯ~�3��pNG�9Κݸ�K�Ĝ��;��R�G9R�@ ��>l����,6Q�Y�d��VAO�f��h@�(�0kHO���X(��~������u�.��������Me�z�%�B���>	&��ű�����0C��^g;x�_��/!ٲuד�f����p޷a�AjӢ�]����G;E4�n\K�:�� ���K�S�C��a�>�ǅ��5�l.ڨ8J �	�m�1G#�\Bf{����G���!�5	7�d��,w�g H[לs���R��R����!�V�9�Y�@x�;�}ƴ|4���Z@�H���2+.�n�M�԰׀ᜩ[0�Ζ�L!-�UK�J���'�g���x&�Ϳy��! ce��,߇s��S�Qw⏴�<8m�5��|E\�����\����Β�.jc�B���׾y��1��,�w5��M��ٛ�rGkltqV0�X�6lф��tvy�Sf�]��n����Ż��h��)��}��+)
<��Q8P�=���,�D@�
a/io|�С�;S� A`ge�IlM����T==G���Ȧ�n{��B;y��-�E0�`�Ca�Ih���}�a�����C���ι�s��6�댹�}��Q	��X����>�
-l#*-*�g�yz3��(���G��cӣ��3�s�H���MU����	��Yb|D�3�H��;�5���ϰ }����(^���DM�
���,��ٟ�.��$�
���/b�Ą���cXV헩��N��ꙭ�6�R�NPy> !��OZfqí�����fX�˚gZ���%�"�� ŗ�j'�<���.n�.e;����W4�'�pc�S���r�"*̶p�E�N\^�/>Yo�-�H��R�O}�V���B��ط9�}�V��ɭ�HY���f^Ι;<�ћ6d��]j�o+V���w��9���+P�>�m������Jr׉����������~��c]Ǒ!��%�-�~Ǧ��V����qd���;�C���g���Y�%���el�,ÆC�~�~�U�Ξ���o�V ��^����=���螞�tߦ��� ˦������a���ƴ�sGJ�<9_��1��{9Y��+�<�c8v!Gh�>�å�#VǞo�v��ƈ���;x/fŮ#�=Ox��vf���g�<�#t�Z��6�B�UJ|5�E��icm�n�AtR�7�|�,�)����
��g�|(����N!��a�A.D\�Ԉyس{�Ĕ^��QQZ�������Nv���抇�I�vC�h��7�\�=��u(��*�6ͬ��w9gE�Q("�H�)�Z`�O����T����y�Ԅ`Æ6�W-���em���[>u~�O�2=��/��$�%@��Cʡ$s�'�D��U��1T��HE����q'T� �h�Vu���8�-���K��%A9˙�pA$���Y]RT0�$�H���걻ﾵ�NT��D�ة�R~=H�bD
'��F�ϴ� C�+T�Y��t;g�W�$��i����@������!�9�u��ǹxhm]�������g�8W����NV�u�;������iG�x���N�B7 �u���7��R�Gl����2뜺�w�|��=)R9���'�`17��dl:�h�<�
Ⱥ��r�D�H����eƘH�Ś��]Z�n
��y�G�Q�LwH���D��\UfS_-=9R���v���q= vS�2Ȣp0�"�`�h6@?x5T�{�z���sXG|�o��`:����V����<�#��&V;��g7�b��QM��!I w��s�|�җ�Y��+hkRbh��ĩ��_#PL��IyF�"j%E�z�.��PI�Ok����*/q�h _+]�1U�$:򀸙�G�0to/|�W�8ԓ��m�jPnΪ"���+W�iAOg>�NB�򫮋���6����Ը_t����l��MB���qjv/�K��]�U
�.
ʲ�Iz/-n�ˎ�dZK5���i�>�s�ؼ�9_��=���Ũ�y��.L��Q�t��17�Ţ5���i��cp���/)Q�N�q�������%���w�L�M�97Wy5�c��n��ȅ��G̎���'�l�	}L����ӿ^�=���O�H�>d�R��U��,PmN~�JsÜ�<��WW�1j5ԥ���!ީ3��9Ns�S�Nw$�����j���֎ķ[M��l7�s�ď�9IΉNX9�<Y���R�j&vc��R����r�\`/F��E���X�m:B��M�ܕ�P����m�Z�u({��Ú��q�\n.�Z*���!q����(���G��[� n̜�	?[z;�a}ʋ9�@��G��X���f�H��n��j>����t���� ��"#3aJ��кK�e5��MR%�[sMWs]�y�L��:�j�;׍�x.�ƅ�Jˍtۗ�~Z�Q�lP�V��pZ����sr#b�آb�Dx���KB��YԄ����B��e҅B��w��Y%[�[��E7�,I�q3�����<���.�䥸IQ�4��؆br�ŭJn-G��Mw�b���H��%F�j��zIq���;�V6\�p5����^�8�Q���GǑ9N|�_g���vnc�)6%��z�g%�u��bđ�T����0ItLT���f���L��]f�>�3�}��F�ʴ����鰹��ID���$#KjT+`�����z�uIQ��������Ç�2��P�t8�"uT\jv�oS���\@�l��輥G]�p�q��\rR*�.&뜛���E�t��V�.�ϛ*����*���k���$rF��8�[n��)�
3�d?�#b���v$�qZ�,���7Uy]F�\��b\qP��s�-F���$1�pE�����M|ђ� ^�z-;H÷t㪗�y��ht�	
)0@>i�A)6�n� G��:�)��eYKk+GE`�ׅ<�s&�F�P�i1C��y*[�i6J�T���X%~'��*��u�+T�����Qb%���w�Z%���*�W��9�#��B�qk2���-ǻ�:<��C=<�ǰ�b/[͸�Q�J[�C��t1�I����U̚�"�r��Z�M�C0.�J���.7c���%�]D���%-�"2��A���C�4U�o���n��^d�n��'�.���x�<S	&��2�A��~��;�&�x��ج��Wr�p���y�[���R�j�����CZIKh�ZrN�]��R��NB�p
̦���	���|���U/�o���xQ���~��*������cI�t�U
Y*��\��Rs2oS��\9�&d�"n����i`����l���^R�������N��s���5�C��%'o�τ�i	w+�W1Kf�.
�O?	� 8c�=Ӿ�=��{��g���l1y&4$�?Ž^�+^�8�X)��<���ݣeW�Ə�=��Wu\1����a�}䬾{�1Z��BȽ�e��	���ZNh���c�}�Bݬu]�"����#ާ�Yd��|X��b[�eV>�����Ͻ��������cTＯ
��DyE	d?����lN���5l=�Θ��[�i��qLul���ĉ�1Q�>����z}�끌�n�A��O���Ӿ�t'}���a-���ryˆ M��Y�dn�M�����SY(�g���Qn�LNyS�am�V]�Km�v�����qӧ�U-m}���~��
p�8ٛm��C�+��S�g���J�ct�m�v�,6�X$m��klf����T#:���v+�	�^��:��u-c.�l�nRҖ�B˥ıeI�A����7h���`��,q���\�8C��N���7eܵ� K�-����3�'�Q�ˮ�P�qۜ[%+c��Wp���[�����˺l����b�n���~|~zs��+�!	��5*�י�T�ds+�0�-���q��ۊ��ۦd�A<dyr��%G�U��	��v�ú1��U��]V�7�]���e&gi��g�ybs�$��vom�༜{3�3#Ee`��"�>����|=�?��w5�5�Ǹ���W�i��=1x{�J�=����ŰL`g��{��ݲ�7�le�oj����n7,�9:Ҭ��VtCc�ȅ+<}e5q���������u�J�����̷2�,ֈ�Yu�5���շ��"�JA[y9�P*��U����c�4���Qjq�����=s�<P�"�wu��@�ia�3H�� ���L�X��{x�[�!�Q���CΆ�DiF��4ݽ��6���9&�m�s�M�oS��/WMŨ��Z�5
�Bq�MB�p�u��]�Ԩ25�OlG�ot���Վn�����y��^WQ�W)*70��ؼ�8�Q��.�+<�R�b:��!��.���Q��:�p�)��M�rCe`�u�Mũ�z�.#P�8�"y���5��\��0C�WՌ�S�'�χ8��P�3���I�����������]�K�w���Go���&�lm�5	�ʁO�	�m%^6ؒ�V0-�9xJ*BQw%<5���\�7 ��Zv�1�W���1YJ����Ŧ�� >��Ўkxz��L�Ѿ؃i���K�Uc�ۻ�<VJ�Wm���v����s�\n.n��Qӓ̒��-Ɩ����qzzk��\���r��q1�����AE��t]o�+����'��-���qj>]q�WT�㈓�9��Y5�˦��I1�>߾�Y�����)�7�9�n���ᚗ�"�> ��eYTBC���!q:�Q|�陼��`�BHkT��J��u���L�I9@\� u#���n-N}�9N$�I������;XW[r���^��s����n�<�޻�af�b8��xp����^����.X���w.�vd�"�Z<*�.��ytơ�T���)��C���n-F���:���Rp�RTn&aq������G�q��q�e@K�\o�o��U�߇*�1���/ ��ˈ�4��e�͕��LGQ;��`K�Ǫ|�'����B.��j�VÕTڊ,'4y���J�,a��X�]�]UL9�Q���ĺ��n&aq���n#q��xl���jy�1D���P�Jq ���n5
��\&+)Q�ҕ�1@:�n-G˥�i�7�I�����x��5ŭʨ\[�+ޒ���]|8F��^v}��I�P�*��NU��Y?�4��&��%̹ސ�m"���nvPy�6|݌:9\/H���=$���WArpi��<q�c�@@,l��!	�"��,`	�,j��"��98�$�K�^���cw��T��ݱkN�+|��qE�Jn-G�19sx���5
��#Q�8�����n�4EB#~�o�f�x" �^g< w�(�?H�T��C�Bj�I��.b�d�=rk�x�2�y˴$�"��\Ĩs�/s�O��b��2݆�m�m~�.ٚ�<�fy��}�g��gnvgi�����V��]]ӎ��1Z�C�?���*���<����t�[-ݔ&$SU
��r� �/7M�:�Y�_���Û�y
�/��p�v�!�D�.7>rd�wW�Px��1Cu�a�q���,�(̨��<9����H�Њb�˵${�Q41�8U��ak4F�F�é���ɉ!QI�BH���P�"HZ<:+`w��l ���y���p��`z�PH��'٫�g��}ۻ�';��k������Tqs��u;�V��悄����yH,e%)���s����F��[��cf�Y]O;�8��.7 ��n.���t��|&:${��.��c��nb�ytơ��b8�ԏ�߭����#*]f��n�nd��-w)�G��k��*q1���s��ļ��ʧ��怳��U�>�?2�CFK7�,��;�Z�39� |�����S�6�3�VJ�v��jk��U���UK]P� ID � a��$ ��&��(R���o�ȃ��%c��*M.��.��|�^����ևC||"7[8/�������L�F�;����^��d38��y���Gi���
�r�L�����xLE�f�������eL����]�8�Z��u|n2��Teh�+8�oWm�4]*J=*狠����7n����<��s۳�u�O��E�T�]vwhU�t�nםx-Ԓ;7q�_$p�!%8�)Ō`���;ڐ�g�K]��j���L��)�kx�@�����S����tQ���� q$�,!�W�~���侖d$b����,��iP�{"��`.O[z��ȃE���!���656���l����:�C%�T�-�)�=�D&e�*���7<Q�-��l㧔~�e_9�*��`"B`�`t�������O��
����m�ry#P��<�d�Ky��9� ��K��({�aϔd\��^xd�6N���$��f<7W��Y�䜅�u�}S)���2O�5W	����=!�*RĨz��_��=��(_�N�����%;é���LQ��Vr���\a��3�0������n���)\�R~R&C��Ȟ[)ԑ��hN���ދy��~��'�|z��x�^��Mpu���y��/�7���5�<��c𜽋�]u���<f����-u����d�2���	GeXv��8�Ԧ	0n�Υlm���AT�h�ȅ)��E�4S��Ou!Zf=��ZG�c�\J��y��{���^$ߪ��x�Nq�!����d��0Fk��=n��5Y��w��ӓu�C�};?�.?0D�~��m�4t�4��C��'u=�]<y�^���omV���Ł�j�p�9���VM8'v�h��4E�ed��yktܻ�K���i�z�Ν���L�q�x8x:B���~ލg�-~���Snp80�{��D���B>g}�;�z̃ᣳ{��~�E%��yr�k�qt��zQ�c+��.���6��{r��^���,�Z��{�L����X��$��? "����r�ǴxdF$y*�xy�K���Kr��t�'�iP������y��+����X3�F��FC*�����{@�A����&��7�q)rGU
���U�?������	�HNǬ{����F�d�Fڽym�{��&��lLei���h�&@)[C`�[�;6��y��VE5���D �n!&)��c|�AC�I��4xFj���Sz7���� HΏW�	�ئ�xb�k�ԯ1�����P囜��w�jy�^Cb�h=�Y��}��|v�}K)u�μ���s|�R��}C$hb��˟k�#\�<�ewrn��r{E8d����\qځk��m�ԗOD�!�m�#nsxu�v�1�,	-�!A+K����6����S&ث��g];�_|:����x�V��뛩���v��fޱ��<��$Ѿ���8��.��xf��h}�߇�^y��<��
����hgF�10Met*|�$wStZy�}�o�����h��;�'4D��8b�B��7b�_��0fg"��H�P�@�(��.�J �x��Mɕ�������U<0 : �F-�y�wZ�^���7�ʤ��?����f�` 
�2�%@���0���A�EZ�򪑋��l���ﺺ�,c��O��\��3������� P�͏��a����;��WB�jήA��\���괊�	��؊�;-���U�J���2��@�zc_*�=����"l��h�����F�'�i���FƸqfƢ�'��J|O��v���{��.�?n(�!O�@�{���D�P�.��a�|ٕ�G�RԻ���3����d�_Cq?/��s?��i-e?��9��n�'7f��p2|��C^+U Q"pF �ʟ��ϕgE}ʓI}�4\A��f�'�iK�f�%(Me��}�!Լ�J|��m�[�h��������+|4x:�d�v/޿���k"]߽�R4Q>���)�i�n�+z��.���R�z��^�M�Ǽ���l���ά��bq�����Tb�	�q��̍�zl�R	I��m��#�BQ���[�t�m�*:;7�ή�ڳ�]��nx�#"��<n�wHSnjQ�YE1�kQX
�UYjp/!Àf��fڸ��24�$Rݹ�U�E�=۳��\��2	�������@�p�ԟsx3�������w���;��c��a����3�ٔ�`�/c�RM�t fL��Y����mW���m5�i�\cGU\�x�$R�q�2�mU�H`F��(rOפԵ�x�9qY��E��B���R��S#l�4�0�Iyy�$y$R_ �-�eg��<�Y0�r	,�����,�+韒���<�L�H�;��g�f���d�6t}�ц~���������	d��!� ����!̦����Ig}��{�����zC3�������6�ؿz�����ē�N���-�cTO�VdE�*�b�8yi���'w�,Mc�������CeQ%&@~'�}�:T�un��6�����*oWd�t#y�����J���]��V�{�fF�Y�]�� �q�H(�I	�ʥQ��2�|T�UX���xX*wC�o��P�S`���c�����;�&��h�z�8sgG�쨝������U�oß|�(��S������o�zx�b� �b�dT�1/�<�2lnp0'm��8{ٳ&�9����ԿV&��5�6����۫0Z�t�T���������Ú9� يdS���a�c���;�S����Biw*<�W�C��6txo��e O	#������|�+U�S9���.��M�љ��9��|1(f[���g�#��Q�[��w�S�1��6v7P��#o[܌��U�бy�B�V���9�;OR��z�M���L�����T��b�]���wD�=���X~�{�>8SO��k7.�>�伱��p���K���M�/h��|Զ��=j
�?G:��p'X�[��v6�l�E�ݕ�h��8�p��-DeS��"�E-�~���Y/��˶0�;NM|�aILX��}���o�L�kf��ʐMpU�3���j��+-ֹ��j�5�5��X�5Z�a,�Fh.u��m��V`�uL�uĳj�m��H�&Y���ޭM�4���7@ۇe�[�[k.�/;�TśڵG:!ܴZ��ݻs�"b��)ܱu�tx�nܫ�m���^�<v-<K'�2�p�4n�(�͠-�a�gsH;�f[��՗B<te��h�IQq�ܝآ��ru�a��k^��3r�m퍘x��Օ�&�f9ɽ�x^��.hǛuy��a�`��^;l���\���	tF)�gs"�ۋ�<skZ ��.�-��%�+T#�G���޾�s���>ڟ��Q�r����~��{wt%܌��S�Vd����D�9�U/���ÍI�. �z�>[Cu����e1k
�1c6v��6�od�G��f3�����%�s�B�yvS��7��<�3���#O�-:��p�=���ܼ�$��'��Y:��a������c�{o*�TE��nLx�g��[�>��yry��&�Ǟ�.�}�Z�{>�^�^0Z)�r�n7Ks�MjU��jL.Q�k���).	�z�3˰�`�9c��v{J���.��%Mmn*><' ��r!Č`���u]������}�V�LBζ�ڥ&�viw��<Mp�I�D�RD	��I'�S�$����1Zj�~� ���/�=+�1�rrV�I�1�/�®�3USc�:��u?{��Z���Xۓf�m���B�vO�R� ;ޗIn����f-�� �;-L}s���"����GG��zC����@�"q��X�b��(���*pKnCP�� �\�:&9��kx�k�ʩ��5�jw2�@��ts��gRӴ���wU2y�\:�&� �mf����i��>x�v�<t�+=o�-I?�G��D�V���S��I<Qj�]��qG)+�D�;�}��A�^(�J$�=T��7�R�U+��h.�"/�� �~�[0��N�у����?Ol�K�չ�L+l6r��{�˒��_|�2Q{�{�zP'����6�{<<!�+��n����+䑓�p{ ��q�|M�5�w���f�N��j�5��F��ə�;AC!�{J����{鼝} ��2*%�~��I�p�';���$�SJ�;�-���f�Ұ���뮱�lo��.C��P�;��%a�c3��ɧ4��Z�u�yAm�UJ��Ň[��~ �t�6QiW�C�L��`�=͝��K�p��v�}"/�6j8w-}�J.{���э ��b�-��ń����%\m�lvx�w�U���x�I�����گSʮ:xA0ų���CF�U��7�R%A%%
��BQ�t���Y�8Z�]�/�p!W��I;��;Q��Q�����׏�f�D)�<��?����b�c�?�Yo��'7U��=�
(�\����{���� G�����h��"��鈗0�Gv�f��߾���K>��'�?co�l`�GzpLh�ܹ�d�I�Á,@[Z��y��}�d��r>n�(�rG}���/�6��-$g|�y��	�)�ܖo���[| ���κ�U�O߻о���.����Do��DIb��M��i�2�Ϟ�i�6w�@� I0 �4w�9'��o|fn-$u
�X����f�6~� �| 1�a�'�rN�{A���Ɯ��iS��Ȫ��'7vn�t��A��	s]3c4" ���6P�S�r���{�o�w�&{[8>{�5���I'-Ͻ#�Y7���Vހ4{��FR����Ԝ��y�v���c=C�܃��2��c��0�q��`�X�Ŷ��h
�6��$�1�_;#W0�\�K R��C׋�EhV� w 3uHxx�P��e�� 	f�?}��R 3�͓��3�����]�W��0t C����/���� �xׅ{�vF����'0�� �t��]�_]�^�q�4n��Á�.L�پ5��FO��`�%��U9n�-�Y���*����k��K��1�GvF1�<��7#�z�4h�D3,���!�$GÑ��@��n��g����f�)n�1�Uɜ��1�/�j��<�R·�K�;���B��\�*�&�[M�Xb�9T��;��@ �+��S��yw!����?J|+��Vf�����I̓ ��� ��� ����b{��ѐs�\R�v]|{j�l�/f0��F��+7�����i�F0�Ѕ�@�B�!������s7U.u��k���Rw����C��}�&�Ҧ/ε�5KT��gz��)̦�/%ܲ�c�4P�<
s1;B#<'=�$���>���M�6L�� !����&A$��eLI�>���TB0ř	Qm��_���#���f�C^����o�' �s1��P���cnq�J�5�m�ùgh'��أ���'+{˗�Դ�"�ϵ_Nr^����NC�=�� ��HG6���	{Z� ��#A}�N����e�j^�2U�Hwg&���/.�GM��{ݛE�H��MoM����{�3h�#����qy��&q��-�p��z�F�'j���7q7!V�孴�l�_Z�ص�z�b̙�V�)�z:�bݪ�I�,���<n�G���y�����r3J�p�|��݈_��3o���H�fp��w�xEߠag�6sՄb��������ѧ��h�򚟵y���}3mW9]P�G/n2���u|_��|�}|rS�^Ѿ�+Ν��k�yq�gXq&6.Y�����k��z���媠�ɋW��͟P	0��^%�.��X�ӌ�Dlد\сYPZv�����)TG�x#o�I�n�}�{�P\����$�E�^ �g��_AnOsg}�  ��S}��Q����+�%����o�T�;�a����ϕ�^��ٿ�'d3=o�{�se�e@
�~�#�N��~YK&I�Əh���'�M��gNd����mS���'!f�ld���3��Ia �������7��i��/���ʩ��ɒ���Й�5�l���ͣq�$��tߐ*G��<gJM	#������)>�y��`�=�4h���������-#:��� O�H�{ې.���S���ْl���Ǎ�=�1��=�jޚ{�5�����G7e��e�z��du�S5���Ѷ���U���q��h�,U>B����vq�ɱ���Z�irFzp<� 'R��vis�5�eb�b7����NϊwM���M忾�ēg|4)�KJ}��W?�9'�����L�e��&��9�g�d�G�� P�C�bp\�߭=�~�^���#���)bK���6�E�OX��}��c��OgS�;)c&A끿LU���l*;7;�{#H��p�(�(����·�������b ~俠���K�N�f{[��{@n�9M����{�G+�˲x@�=�S �������)��[�뫢\���[N����L(�]�NA�䣚���$��J�"`��X#�����)هgf��1��2��Q!!&`V!Z`Z�w2�&��������˰~�M�G�o _4L�w5�)�;�`�j]�:�kY|ロ:���ityM���B2M��Wp�%p�ç.{�0�I���$�{����x`}
R䟷"�GD���ټ�����RKy���Θg�X��m4��4���e�jA9�nL�\Aİ�m��(�̥�+nTη^ߪ<�yJ��Ҹ-�'u��ĥ,I�����Wd@&��&kf��nY�܈ĉG�s.��|Z2mw�. �M)�HO�Ib�F�K�r:ʧM�HG��1�0[n^��vA�y�<�dc��t�1fѹ���ˊ���6x�B%����n[�]��� �3��d�;��ӻ��kM(�-6 �ܽn����j�nPF����-�'����lrD��T4���3@�AX���I�	Q�L�v�������[{տT�N���_f�CF�6V-�'�pL�l��	ho��[f�|0�m����F�����w�sTz-b�r��VK���Y�400�i0m�����e�!8�5NǴK�,��_}΄��4�&|!�eg7�'��{�2I,�����ڄ�^t�u:h�i.T	h#��}J���x� ��D���JT� ����d����;4�1V�"�d>\n}أW��A�N /B��9�8}�R�g��Ȁr�}�7�,��Yjyl��v��v�B-\�i�`�wv�u��K�^�;�%�}��pn�-���}���Ff9!���7��������g�TL:�U̠�f���Uy,_��;�����{ʋ;-�F�'���`7�(���1
�P���� =�0v�8����R}�@;o���`���n>�� b�ڞJ�Ɉ�{�`�FP��a���׸�������{�+,���0�h�o#Zch���]DPzW�US�"�x�0'�!��h�>���\�O+��ؠ�¨ꚓV&q��R��[������lz�ӷ��~����?Q9��L/�n�]�b{���㹩t�z.�= �s� o5y�"���{IK9졥�ڥSĺx\u��^�Y�g�����OE������{B�E��y�\}WA���~�/�����w���,Lث��J�) ñ�)%�?�v�W�Ѣ�'�t=�s<�@�Wm�y��ri�LlӱҘ�ON	U�)ն4pK>�e�yu�m3ծ�Imx�j�������f8yz��no8&��ώ+l�!ͧ3���V8�(q4׷�ݷ���#�i8��a	�m��[�w<�޶	<-=�;۷6ݶ2g%�����k5��d�#�.��TU�Q�x���6�I�:�v؋0V.Տ�R�!,գ[��g��ס�u�]�[9v[��%�T��;����hl�I찾]�J�f[۠˘�6���m� � �- c��H�ן�Ǡ�\�mPF��uo1s2��c�����|�ou����/�
k)ẁ;F�DĠ�$���{}�i�\�ÿ!�B�'�<���ju�	"��%.��"���1xůz��v���� �^B�~G���n�E�o�����6z�柢�|X�
��u���2�yA�D�ظ�l��"��e�2]n �G�{%�a�B2v���K�dy��3'nv�`���+di�X2�9��;~���ޱ�mPְخ��"P���Ґ(�*۪9�u�]c�v�a2�s&1׌�̛$�Z^�ٍ.%���N�XUN�ju{�z���JVe��b�Mm����z߾_�B4Q��hO�%$����^���5/��d��KzQ�r�8L��ܨ�ku
�R�g�p�#1P�#�K.+4�k/5�Աf��g��g�x<�Kvz��ܓeMѺ7R4�q�]�k�����BY�pT�C�Dlq�$o��9%̹8���N!\�s-�~6C{��
�D�Pp5+qg���=�o��֕�ˈҺ]e.���*��&e^�ąs�F��\��ou� ,IĄ�D%�Ƥ�U7��	���09z���^S�4@H^<k'���'[n'�O=���1�(3�'�p�Q�V!��Q�T��)t�[[���7m6o@f���f
2���Q(� ��}͓&�]�a�FG$YV<�։����f�c� �(�[݋�p}+��ۗ9]���������c�<O�����0Rfo!f2m#�%�<�/�N��DB�`'	�ˠq!����X|��UO��e��y���2Q��n��4��eVG��n��\�.c=��- L �dƮ\JI³�q͓�튚�s�������i�o�h�O�~Qe��r��mz�ǵ��鱻R��;�l��#g=S�c��g�f�^;:w3Ů$8�`�Ų�Xm��7�ߐ�ϖ��md�c�{�w4�U��u!��G5�۝����9�^�"�y�I��h�'���64���zݳ��i��`0IeG����7��g-��2Q�n��g2�!��	�a���0MÁ�8Q��� 'R�S�I6v��Y��/�F̺ʽ����/��x*@m�J���߶���JM�O��t���&J;}M9mM�a#�@�TV�5Й��RC;͂g�!�w]m�306�0�rjb�}R`���ã���:��	��(Oq1e��n�خ���������xw�KUQX�`5�z�d������E�zf����ٴ��>�ˮT���Z�.��s:�/���m�˛�ҵ�[ݵ�4 6�q���� ���?W�H̑�����g��/K�`�Bud+���pSFn�����6����;zN�3[/r'k(XhLLL�ai�:٣]}HR>ɧ7<��O���p�-f��J!#Y��g=�x��>�У`Jʢ}��kx8R0�7�?3��� {���^���Q\��Q�/�n�~썦b�I���ޞ��;b�z\�]�>�t�G�`��ݔ��OO4�ns8�lF�h[�kr��8�j��.����$������G�;;�����S��8��&ux�{�S�m�ۖUouB���L�!�]���Tr4�	�X��Zh�L������'t��� �vC1��F{�J��Lw+�Cz�Kl"""8�6���m�����N��HSx��+m���k��e�����������օw�(dM4ƚ`	���Vf�-n��A��c13�)׽�A�C�`�C=�ײ�����\0L&Yk�8a�K�A0�D��ą������vDy#Ύ��-#ت��'z�)���*0�T#b涚���1�[�t��:GowGj�u:�S.'/6�9[�&`U�oY����+��
��aL=������uѳ�~\��:!m(��b�og��~�<�yܧreZ=�L�y>C	����H���fٺ�}�0�Q�C�:y�9buf*/n���<��nXY�����T��k�g��N�	[��ݧ��ػ ԣI�<��t�P�Lű�˷2�Y먾�-�:&,T	aE�e��h�0�P����L��{X����2E�}�(�7��V
G��d3���_d�Y�>#ޕ�n�̜�	��X7;����Ѐ�B�������yװ��\�{�<��{)�/&�"j�\�[���M�gvRw���o��X��T������-�_,����}�2k�����=�`+����	C9��R;�17��>i^'�{��^0-���/t��r��o�=|7g���~�����
��[ǀ���NT��
~8DRD��G�T����9��)4���_~�����-�B_LL����˽��g��Bg�7�2GJ -��U�f{���㖛��,��]t8��%eQǪc�a�]y�	�M�P����'LM���gigvkoK��N�
G%���� �(�m&{�<b������:<n���)��/�i���d}w?|k ���&1A�|�iq�dg!ǅ��=�6��R��{�swg+�j��W��3s�Ft�V���h�l4TA �2���@��s�V0� 쯬�/���O��l��]fWLUGh+�3]P#fv��3�EE�v�_������88K��Sj�ҡ-����/m��%�r�F���讛��#�%[7��*=/�����D>S�U�1�}�ndo���t��n5 X3Mu�B�s/�������5#d]����h��3�;�����b0C�Ak
�D���)Pm.!���Mt ֐�x�!��"��3`B%=S዇*)P~�Y$;=��N���{�a(�͌7.�5��2�p]n*,灼Tgy���Y�-A<���Y����*K��M��U���*��3Y��B�����E��%1��6&1��J�92�u��5�r�ׄ!U=��t{)�!O��v?� %�L6�6f�H�������0��4
�7�zV��C�R4P�BM��.ȡ�8QS~��1.��k:	���3}�`��}���xē�R9���\�H�,�:P�S�9A#c��rF�1�3h��Z�����>�G�Og�U��x w+�0<v��xԍ1
���R�$˥߽��R 8j5\Y��4xU>�����	t!��u�u��xr9}��Κ{jqR�U����4�{b�
��%���='q�,�O�{](�v�Μ���`�ͱ�E�WM��ך�X�,d�N�q��jء�cR}��@�	@bq	7<���s�����TOsi=ȫ��tJ\݁�+���	:�Y�tb� wf���l8�N��HFD�g�sk�4��ԑ�Qj���|~���Ps
C������������g'��It�F�	� �A0�@"BP��7=�d�+w����G�s� ei����h��� ���VZ�S��U>x�O7�K��y�"��h��@���He�0�<�x;��o]W^F;���D����)VF�UR���,��z����잲)i�nV�<ʹŏ��DG�%���xMM@��*j���M�>����H��RE�� �&�����TX�dY���M��s�:u֨�0��b9gE&#F���KɌ1crv"F�`��'!"1_���ާd�ΟI��ԓ�����mq)ql��,�P�m��G��A��s����]	�^Op�H��Nϲ��J����g�{�K�:��{B�i�\@ӗ�S��v��D��zb�r��MI�36l��\v��Dp��ݪ��Ǖ%�v�	jC.�/��c�d����Ƕ�e�� p1u��ӳ���O�)c�ݺ"�]?MF\�"���u��ހ�?c����[9*/s/7-^U���%�t��w*��*xw�i1N���sWzR���L�5��W���k�}=-q嚽wN��$�4��;SP���&�b۰�����=בwr��_e���
�'q���˱|��MkQu�Ŷ�E�wiݤ�^�-FXa'G��ym��l�iSsl���L5�Vj��nXK4�<�ѧ�u�;��[�����t`�qnC�#�6��etf1v[��%�+���؜3x�-�V�(�i^mK:�ln��Z���Լ6K���M,�J�58�4�A�܀�1t�8����h��KP�s��/R����h3�qDg��g���K+����+�}���/��8�8wT�h���P�uq�Lm��;���9u-�t�˭\��u�����WnѱS�cm��t����
nw�HU"��6���/���w�3�]E5H�Ryj�w t�0D��1�U���w�����x�{@��:��j�
�U�{aNI�*�PRou�N��oJ:�'�e`֛�l�}s����w����
<����H�{�[��>Y7����s|Hdh�)���v�}���(w���kH��/�����/#����rV��ɋ�5�J^�sy�
˪zDѹ"\�ruMMMߥ�����tEO�7�A)#�x�Bc'H���6���Pќ��O1�a���k^�R9J�v�`�Ҥ5��`�55864�e�s�N��I��d"q��I����K��6�5�,�]w����A����}lu+���Y`/M���	~=�Y�g��6�S��w|�:{�;^���xi�n�`ɬ2`�a�!��	|��Uu�W:tt^�r�#ù��H��#�W�K�[� ��(��/��c;AT��C.�%w���}<������x�)��f�z<�����6]1p�c�MorȂ;�<��M��`;:B,x��1L��K(��f"!�ȬoD�ѻ�wh^>���V�KYW�*�V�A�"�/:F�v�$�28��=��1��xt�:d
灺@A�$�-�0 �a6a"4�9��B���{}�d2.<�
��7��X񛥚9���p�Go
!��;�t��M�t�tҭK�Ԙ�5�����!�&1Cȡ�D�Q�	�+m?y�"��$��J�.���u�;O������/d��K#H�S5�dN����l,�<D�>1��j�p#<%G���0��ǗTWdJG�{&&�1ZY臵�g�[����}\�xsǙ���'�k��]IՓ9�6n���p�k�P�z���M�%��٦�g��)�F1�M��N�Ã�,�]�T��71Bk.�X�h�;�A��49�M�Io�V���^�&�5G�_S7�t�ˌ�`�AOА|l��,Ǆ����[��b\K ��qAh�|C=�k�G��#�l̅)N|��Q��*Dl̫��:{y�O�B{�e"1	V�U8�<��^�7�G
S���őg�ZR</
��x5���<���Acw��56�L0�&
h�A��+�� ��7��@��7�P�_X2�7�#�*�Y�G�n��=}1q]��F�5X����%�L��4�W��T�9AB�OO)�R�i<;���|5P�d�d�6�����8>��n-e���UuCu>~1���)�j�	�$܀�GP��Y~q�U�yӰl��,�����AvO"��!�w:�љ�a�Hm�JMJ4�h"G�5�)v���Az�_��W,Ų��Ļl6m�q ��GX�ft�J�дy�):p���H�#M{5�/�����}򢟅�t��if��bM���M���f�|���ӛӤ\�1oQ,6d��ܹ���Z�&�L�|���yγ[v��ZΗ�ײQ�T��^m{/��sd�q���å�a���yc�>[y�V��Ƨ/��'���1����pR@� ��ڡG�F�:��_(N1V��"�9ܪ��1Jǻ�����e��` l��ə�C}�\�$�Ϗɶ�
e��2���C9���7������|"�������u��%Rټ�*[sHu�	���z �d[U"�Kۊ.:&#3�Y�)9�)X�f�t�NldI`z��*�SLQ=P�~3�����j�hͳ�s5m���|�?�~}:.��� ��0G��4[�|��pD�M��-mL����W8��]�%7�w����l����y{8K�1�3�e@=<a������8\#o�ԪZT;f���ԡH�rĲ�o5���3�%��q̫�3ۛ	T&�^;Q�W�l�����1�6��7��?e�N�6�yo9{��In����M�Hr�1�7=��fC$��i|v���Y����j�0��(8��a\la;ü��k��w�|����w����	����> �b���V[���v����"�36p^:����46�_W�9CM�?ikU����&�R���ʺ�õ��Vd��7�}w��i!-Ͻ�z��|�؀:�\=�ĺ�̈����}�ϩ����<½7!㱦���>O�������x@ZdkBL��f��q=)�Y�QѸk��0�6Ա1PQM�a�z	ٰk-�wRQ��e�o�^G����o����{��c��m�Wh$����#$�jUų��\�D��L���m�d0�a�e��!:��&���6}�chp���q-yApQ!w>�^Ew%K��j!6���\��:�Z�T����2,�UKj��Z�8�r��ی���@�����fL��aLv�����a]	�����U��%�E�j�B����,8'U`!�/�2���z��w<h�q�X�)6%�h\��o��9;�'��V��!u^* ��x'�Rs���/�G�Cٮ�2˭c��dg�7��m�ΑhF֪�[�lW8�\�z���>�>[�ZX�Y�;����7.�Ռy���>��i��sOM�w%���X�x��M-3@�(�l^fy֕ED�e#ZE��aþ�}�����طm����șv�b=����.�S�|�H
()�	���,��2Q^�kt���4�h/Z�9|��>!����t�X�f�s��<�=_a�W�;.r��S0�ը$YG����6���$v�K�Y7�H�i(�T��I$2��UW��iw�t}�~o(�}'U�/M)�z�i� �_���ʮ O�B�F�}�u/�P�R�.�����a�0w�3;�-�u�g�ժ�կ��U�*+��eg�Ǒ����IK-B J�+�w��_���`��h��@^>	pDDB��Z��I$������8�N�c*��]ys��W^�tGt%@`��H����za��_5�vgN1KL�!��p\A�ĂQ��RX���`���`�k�����s����D(䖣�ƅ6�PL%�s�z�l�4
����':������h{z�@�����׃���p�?k��u#Yd]V���WB.Oo{�y�ާf<��3���5Ҳ�gViv��`����X$&6�g�6z�۝�6�5j4j�سj3K ��h�U�,لC�_%9S��-A$I�M��D]�}P)\���D�q�Y]1�өi�/�F�2iQ�T"�m3��Wf�+��q� ��q�2���%��se��v���H�r�"a�E�W<��Jx8���U�jz��TWU[�s%�9�
����@]hUX ��%�5n'�Y�N��P�B��0����^�ӟ.#!9��o��'���=���|+���E��:T9i��'y�'���JO;g�f|hm&�F�N�viСt�A��o�C��P��I���`� �ZGĐ�h���j�˰Oxf��O�r�k�F`m\n�ь%k���%��Be���-��U.��6�VD}*�hW+�� ���Q^F�B�3�������Y��+���ɻ��:�.z�1�]!� ��_0:��$H#�1�@E��&5Y*�V������_�	E50�k�v�-�mN������N��^^{�ޞ�
фT_�nUpRx"��r� ��=V
��C����n?�_g���K�/���P�  B��R@�E�" ��'�4�hv����X�)��ݙ�O�ë�2@o��ABAD�Q$A�YDd�A�H�dAEVDB0dUH@T	Yd1�����1E�� ����T�8����k���TsdUD�I	$ �@XF@A@$Q���
�
�u,  �@C1QJ�! � � ��� �cA$E,��@
)��3e!.�E)���A��>A,�!�x}�?I	@!0?��?̯��*���o�O>�y�d�E_'��~?���=P}1}Z��/�b��}��>+�����֑����'����V�Gä�>��'�o�z
�({�#�W�>�������E P�DC���������>����ч�
�o�� ����'�!�?1>�O�DC�'���~�|��}��G������d�T?C�?�~']ပIYκ΢�������Q�_˿����
HA"�"�$"�"�* 	"�H���HHF H�0�b$X D�0�$"*H @ 	(H�B� �
@H�B`���b��$B�b���H@�A@$Db	�$EH @"�
� 	�$ �H(@��X�A�@H+
D`	�$ �`,P ���D`	�$T�$V@ D�@`	"  ��0A�Ab,B  �H���F ���D��H�B �3�D�$�E"P@�"(%
uy�P(�����m�(Pg�i���������a�>x{C_�k�~�'�}|�������r8���Ǡ�� A�� 
z�H��>Y�1�a�l `=��>)�'��{����#�ޖ0X�l$��'�:��_���" ��l������=�ս����F!�}�C��� 
���H���l�����vh> ���G!��8�aH�
��211�B�;A���G���2�췻i�
?���d;�� u�F.� 
�ޏ�����P�w�DC�_��=H{F����c�����}1����g�C������c��@O�G�����v� �;��}��|�@=���d�gG}�>��:F��ե���>0>C����z�ޛ���W��g��v���(d��y�b�jC��=>��}nF��@��=�t��ES�&l��9Fx~��*������P�����; ���2��{���@=��R��~f�?�/�z��A�z�!��?5����p`&}?y�<�.�p�!�$U"