BZh91AY&SY&���_�py����������a,�0  (  
         P(    �z)J"���D	T�TB(��D�"�J�UIIP��J�Ug �R� PP�  P
 $ @
�� ��-�"B$���Q*w��=�=L�^�=n+�p��ld�h��w��=TB�
k��i��99�]�<��W��!����o6�p�Q����.�9��̫��gS>��_|�*IDUq@��!7�8i��z��Ӯf::���wg'�{�W���@�>��� �9)Q%QI[a}��n�N	 ��3RX(�P��1Ԅ@wP��w`(th2݀����N�}�z�`�
8 PQB���@���^�z��@נ.����tzhꈥ�Q$�JB���
"ܠ�G��Ѡ�vj�n=�=��[��VgF�zJ
H���ǽ��=s�ۄ�7`�m�6�z��M����UDH7v0�+�/\��΃^���a'CCF�Zo
��-���T �'W�}۠#��F�\�C-�[���a;����| :     (   �~ �J220����20��#!����JT�h�`!��F&�2a��U$ѪQ�2�4db  ����I�#@��4b� &� ��T`   	�0 D�F�&� @�4�#HH�h���<�=���=^�{8������~aPT�UA� �S��@,F?��� ��͊�H�A�@E �D�7�U(O�  lD��A)�
(�E�?g�����v�Pȱ��.-�������;'ѫ��'��~w��dC9�q����r[5�MN[���76K�:4�����2����K���WB�X��ԃ⬰����&�eD�GF�*���#�s�	�#g#Yt��'N�!8ӧI�:�,j��[��h���4O73�E���;���nN���ۈ�]�F:��t'1�)��1�d�;1l���ًd���;yM�w'��&1~�
�{H���!��ɻ��Yv��J�Տ�D������B� �&�	�Յ�#��q�7�8�o5�e��,xKm�$�|y`�D�9����:j˝���3;E�R\��1����9��B��o$y�B�4�d3��Ǔ(��&wW"c�惯��Ev��s��z�4Q510\8"]�F������صS���G7(��Ok�!��Kͻyb�"9dXcw��-�#�u+����n����=�b�e�gp����N՗x t����݂5�Q�#���n�C��~
��'P�&4�f]d�_D�o����Y��� R[I��܆oώ�<y�mIH�4E�d4��ר�k�1n7ðhV�b���[ǎ��%��R0�e��<rܛ����NA���' "�`���k�%˳��i�"=�to[�KN�ܚ�g��(�s��m*�pK��gp�f�[�dr�\��V!�m �7VO�To36�ʠ�"��ɵA�"�T�T�h�ۺ5�̺O.A��p���ǧ�{7���mVe��j34F�sTLs�'�
����w���"\�=��\p���'Ǌ�⢱�+�;q�ٽ[�N���}�n�/&:`պ���B]�<WXv&z���]��f�7��)�(Dx����n�\yf�)ew�b��	�賊4|/�F�-.��
��=��r"&te}V�y��:�9�h��qD�n�:�1i�G$��p���f�]�^�y����'rh��݃V� n)��҅�Ӱ�iGT�a,��=�ugo&�n��u���o޼�V��F]QO��ds �P�.��H-q�xY�G��q2zD�)���ؗF�]Hu�ݚlv�os�ί�Ҥɏ\7..�E�Y��%���vq�Ց�U|r�a@"R�ʙ�TÄ��C�������goH��ϥF�<�f���WJ��`G@	}xon���J�����V��HD�q�.�wA6ޙ�%�lt78�ڠv���ވ�:7��aی9���ۣ�k:�ցza庖=е��s�η$G;�F��]�x�Uκ��Wl�hH��b �u
�Y��U�:oLr;���H�E��s�Q�\��{M�oGP��&uM��wsJ��ZReni
X�+^����٧��;��x_Eذ3��A�3���%�MYgb�y�h���O���˹hT%�i�*�Y彐IT�T�.%/t��`7T���]�Y�C�z��Ǽ�.=�gmŢ"x��!���|k�� �$��r.J���X��r�Z��[�����H���:��k4��7��|�ӻ_7N)j'w^�
�E�S8��a�b��{rگGB��Բqx�f�٣�0T/����Eⴰf�ķ
����2vnAp(��BM7���h�`\f����=:z��b�{�f��� (�.��s[�Hgb���j���nt�i�.r9��Tܿo4�[qi�)g][�T���ܖ�<�Oc�ǧj�u��D���ܦ�9��7�͝���`b�V��8]���w�D�N�O[�M�]&��W8)-�n���I� xۨ��p����O7������j;�����iG��Ǜ����|e5]���~�ӝ�0�=Oˍ5�2�un���v�)��ӎcs�X�xT����i:��p��X7zu�K�7��Fd���fo%�@�"ߦ=�9W� �aG7lG�n�w�6�4��6t�|��gc�KFۜ�I���XVg�݇q���#뜔zY�8<����=O�����=k
SJ��X�wr�XX(p������`��n�^���ѥDp�wront���G�]�ݻOou;W��gB�S]/=	���'\���X��GtEr�m1���1�X���CN���hPUӵ�1���ˋ��O-Θ��xK�-�9pH���G�dx�n���h<��	:�b:�=
�7I�:Mŉd9�.��9��.�N	3u��m�k%���&�2B��c,�������~���L��sz:�0�H�o�8���ͨ�IN��e����F�{y���]c��qg^K��0�>� ���՜�t�OuP�11$����rmOpW��	�$E�� ;��v����@��s.�E��2��8�7�Cl�C0��-vI1=����˞@1��=�;	��N��� �d(�m���1p�����	yɍv�aK�P�;yU.MO7��9��l���ֺ���0i%(��(ؤh���%�Xd^^t�D}��⺷�*uh���%��8>u4k{[snbޖ::e38tQ�<c�d͢�͸2��C��Y�f�+8��X'A�d^a�Gs`����78��g6jD�f����n��\������٤Y�ST������ZV��^�����g2��TX�w��+�83{e�}���83�	H���&Z��3C;jn�qKB�Y�V�F*���l��س�șe�����û��ܒ�Ɛi�]��{�F�ƍ�RH̷�(�dEJ���-�bö�׉���ز�sF�C|�l0�t[;����ˁ.��t�
}AN�������s������p+"����Ϣ޶>b�ӭ0Oj�ga��l
��eŢ�:cf��	=�B�c����$�	�m����L����Tf�[��Iİ��W��Q0㈷*��؄X,�	{{.@tH��jի�ޣ �F߯]y�`�:��雓��~zfrM�Ć.��ar!hW8k��,ރ>�A�nu8������c&l�}�o;�GI�;�x��¸>

�0L���(����N��R�ÁN�WL��kp����&P����g.�qX����.��"È7�EV�2!t����@'<�Jnmti̙�z¨A�.I�n�ֱd��#�ɥ�빷�G&���V7���l� �NΫ"×T�Gcpk��U!X����T1�H��Lv�g���|��b�BXV��e��Qz�u"���5�*�5��VE$Y���L��i��ꨑ���l[����]�I���R<6��dm"����53_'8\*��JN4b(t�N<(W��.��8�U�dJ�4p�y�b:�}���c�B�Wp�]{���m�ɂ{K�Ҹ���M(-8�]ɫ^.�^�e�#�g[x��Wwh=D׌�S�v���NV�Y�=�9�5�Ou�1����&E���
�!6#�%G� �/���� �"3Yj��'��+S�X�s�W�F󎩉�=:��P��4�'7�����x��[+!�u+ql�m=H��)���	����Q�=Ag w�3h"��r�\^�;�\���FuJ	S���Z� ṅy�9eL�-���s�0�����L,�Vj�p�+U��r>|vRA�w&,b��sTuݘ�̹��>�8��<��๬��XO3U�X�)+ǲϔOr2˒	������-l���oj�Ѡ���fǸ2��.
gLM�N��n�}:�[�6>���Ѐ��`=�Q��itT��N�Í��,v�LFW�+�����F��0�r C�L��S��c�p{?�q!���T�g��'ꏗ�#g���^^���Q�4��~����Sy=�=|��tx�P�tJ�T;6YR�9l.Ч/b��Q1eY��+��22��4���0��,Њ�[m7m��֓�.(�V
������!��ؙ�G!�j�5��]XWcV�@���[bEc����ķ5l�4¬�����]��k.�Du�i�(���fGYu�Ș��y��%Eغi������D����nr�@Ж$0�Sd5b�lr��2�v��),.���{�;�����a���K&2Y��[49sש)Z]��)*�k�eil3)ĺ����4�A"�叐�6���:İ��U�� �T �5��S�jU�X�G�����,ڕ�e.�"V���ƀ@�Fݭ#5jK:�q�Vd��+,I�A���P7cXiI�;�L��su6����R�!�M6���T��T���a@m&[>�{{�	��E��[p�ѳ-ҙՠVV,4s�3��`�"S��f�舱��Â&6bQ�yc�`+Df��頱u�PL$sF�iI`��X��V.Gm���Yn�586�Qp)M�Z�i���F�k�iͺQ��h�m�I[h�Յ#n��v*n�42��pB8��
d�ڷ�g=B5��\�;mb�H]���V��2��&�RU2h2�.�E��ErE�mٔDJ<���k�����8>f������^�c k"6����m�Ye��+ǯrЄ/
V����
8hJ�gl��ñ!���j*������*.��Fl�V�Ƀ7S-�5����cq5 "ܰp�J�Y]6b�YMR10�1-�+�i�<'���,��[5˳7���714��iF&E�=��|�Z��[5��f:0�;]��4q0mnMm���!ɦp��c�7**�M*��W�۳ej��jd���"�؎K��mH��XA��5.�3L3X�l��j(���)(B�KEe[�����i��)h�Ђ�ڜvP���DƭİS5t�RƔm����\�E���+��A�hp%TlL�4a�it�խ�p�0XRn,����,ͅn�Em�*�Yk@֦�QT�lk���d����I��-�� ���/B�f��]�q��t�H	%ҕ����������Ж����FW1���`Քe�65�l粰��\3ku1�E�.s�;H�cm)t4n���t�y�tn���F%�������"�sx���Y��s�F^��C!���([-�b꙳3,�n�h�1 �sr[���]��w�M���"F�Te*9��`p�6R$���(�]B��)%�[���3������@]���mn�f�A��11�4��U�GAЄ�6h�6����n��hZ�R�&
�:���+p9�l̀�IW^Z.PL��136�6�uH��k���Xc��9
�6�\�H��XXͮ9��d��f�Z�b��u�Lݥ]eU���������sHmF��)(���"�̸P�҅0v��a��X��"�C�ʓS!���3��ɥ�!D��J�8�7/�V��#�ыY�Ǝ(C#��A�J.�B�4�u��mn��J�"@�R�Kv5!��n��ɹDغܬ�Js3#KNh�CMu� �KX<�)��l�!)�n�&WF�c1���{EE�:���Q�8F6%��vC�#���E4�֤n�X#�nV�jd��cvE����U�Yh��iMhVk,�P�n��m���7�l�30�ۙ����P����ٍKP�"��jGsE�v�s��;S!pZTuĸ�a�0��E�h\�+b��l(����-KQ%��xMB�\�Rܑ�1I��(�,5(]
e��SQ�)b� � n��Tm53s�n�����3ZPJi��-m΄���ծ^$XE%���U��h�ٵ5ڍ�0%���J�JC፲�a�Gv��!��l���0����km�㍫+%�1]��[Zg)��)�UmGm����M����]�i�����
If�5��IL��&��m�%�B��$��*��R�KC�X��i�A	�ЮŤ�[��"a��ba0�1�+�4beu[�a�5X:ڈ����6��ɘ��Z��3��n˜��K�/S�vc��lcai˯�[�X�s��b����V׭�f����Ρ�Q؁��6�]X�0MZ�͛�#l`S!��"Ǭ�25��uЖh�e9�MÅڄ��5�鐁K���"b���ܙeŖ��&eIH�)JX�V�a��F�bs�ef�&"�j}���ԉ27����j�zחo�lC2�7k�K&b�L��9f�̚�I4k.*6"�0�]�H*����en�4/\V�W�7!�]�뜒�1�m�e�.ҡ����zE��ٱ�4�4/uv�u!��F�ᆴ\�Z�� gBR\��:�ئU��Y�q�꽶KI�[t����`���֬14K�c�\��l���C]5P��굍$�J0�̫bR�f��n��X�0q��bHcD���ӂ� �\�i`�[[-��R��Q���tR��
�Jͥ�mqΡ�1u�V�D.I�2ڏ\kUY��C��Őn�ِ �a����I�	����͈8�8tH�2�,�cv�h��Ԭ�ba��4-q7
��!��3���2��VWu����#l�v�����(��p�1+�ܐ�%r����;U�g�2�V��h��=,�e��(�4�1z��Йۨl���)Qۂk4yC�n���PV�����ɝZ�W#VU��J�[���kp4����1�\5M��\�����\jl��%��î�u8�`&�4I��˭� �E��Pt�C~��h����DP��,E@&��Ȉ{�O�/���~>�Wg��}g���'<���s�q�Ǩے����u[p�e�N]yo�����𛋜$�;�Դ��_
�������}q#sW�°�o�N�+M܄��m~ʼ��<=��/-�뽝�V9?��~��{b�~=��d��zya�
z�J��6�,���$�*�����i�v%0m���<E��7�rE��b��Gd;�r�wOV���Z��ӓ����;�e����i��Zn=�(�y��c�p�Tc{�rS�+�>��e7޺d�^E�vt�X@��-�=_,{ϋ�$ջ��b��{ƪ�k�^��y���:Ѓ�p3���r��]���&o2���徖�w�4���~�O��އ1kL���uzYf9�{��	�)�K&�t�r쯇�h��I�3|��&�A�`�˕�|;г�:���G��޴1ː�ٽ��o�y{����z5�t/'�uB�ݖ���d8�}�;��N��sY�l-�x�Fz��v �Ks8���᳚P�2�
t���F�i��W�]�琝�G�0�Ò�4�3}�e����]�	�`%�VI�Y�ytڑM�� �ѻ?c(P͔�vRj�Τ	J\s����:���2������i'������3�-�׶�כ�����8�ɶ^K����o4Wv^!�\:�� l�3�dW�,�]��6��=�FÒY��zo��&�{���{��r�y<��uJ�Ҽ����w��Nm�� ��
ɏz���Z9nA�%r��/�Wsʫ�q-��A�������F$G�q�eC���4�^O�g����È��w#��՜��"^��_�!�����r1��@K���d~_K{í��۹�-��:�R<��V?`����X;����p�V��h]�hr��p3J)U__^$ίz9�U��q{��x^�F�v�ӽ�R[�D�|�`M�$�橥;&n��3t5��mk��y��Y�N��M�g{rzu��X��T]�?{��I�D����'��B~�m��&P.�zBX����q�h��c�xr�{����D)ACj�_z�z�u{d�|$}ޥN���DQ닍KwyǬ���ˁ������G��dx@l��/=(��EΑo���x(]��K�Ht5�����R�t�*l\W���i2ֹxĭ=�
�Y����q���(����z==�u/4]�c9��-K���k�ѧŀ�\^E�/7�Zu橍�[�TŽ��b��7^���� � �h�y",[��{}��41F�5��O�܏��w���~��r��C=�S;�5{=�=Ç�o����x}��-3{7�'l���9���YZ~��!H���z] �N��?s���2��i|q������'�݋yn�%�_�#cI�P�7�.��VKa[�5�alU���{�w�=�`ڻ��zx_v��*)F�j*������z3Y�^Ɲ�k�8GϢo�=O���;E��6���x��Kس��<8%�_o7`�l��Y�]�oH�0L�R� ���y��8N�}����Y�yt��]�����'�Q��g�'݆!���P;�6�u�k��'����o��{��ݙ}���Ü�ȉ��Or����c��i�hs����v�ur�ن�4_4��ga���+������"�㋚�(}l4�X�������%�Q��<�r"��G���c�|���z)�{��pD)��%�)͚����ﲔ�dњ!'��ߖ�W˷��}�]���{�e1�7L���E|�����c4��T��`�x�{40�N��6�.�r�C��H���9��gg��M�tŞ����f����4q��?G�+��w�:̽<�e�;��oy��I˛��5e�s��r��̽�+��6U�Ayݗǖ#.��}�i(�goR"q���p<����8��{;�2���� ��D+޹�v�r�ƲSWV�O<��|�˙ȡ�,�k�4���CX	�K(��5��T�
!�3�L����R�f�=0�/�?9���y<�y,��1�xn��~=N�v�"�v-G�z�l��z���ưs��#x|������>5�W1k��g��[�=��~W�P�y�����6���;����_v�>:VCh�;:��J�'å"if`��!��:6Ã+6��W�^&���fj̩݃��v�1�#lVL;u�����3��Q�7[�it �)���imn�����j���lܩ�x��&w�c��v���=y��\����!�5O8��(���ݻ�T*7
���ϫ4x+7ԲVť{k2���n\+�RL6M9��������]�����.��m��l�=Gѩ�hn��$��z�+��;.��ۚ��\��H�n��&��_C̝" h;��I��x��:��������L��[v1���q�[��Hӟ!�3oj���þ����Ob���-=Ca@��{ޝ�^��w��{s�������<QFlh��Z�e���f��ۨ,�������c�����O-�oz[�ٳu�����W��"����N/h���f�mu�-��'Bђ���èh�%�Y��ɶv,^G�/�ޝY �����e�r�����=�͘�^�x����m]�W���*�OY�W4�ya��Y�G��ϥ�a��>��@}H���ـǝ��ߧ��9.oȕ�_#�AL{G{���}z��}^�����r�^ɫZ��w.��tu �d���G�e���>����_-��}�S��i=�ʄ�wG˗��ǆ�x����Ի�7�����K��ǞǞc��x�ç˒ӂ�۲��=T�5�]��!Fj����i��G/�Ȱ=��6m����Wk���d�yWۭ�s޺;�(w����]����15������Jҳ֡������홴e�]���v�F^��wެ^�#����q����ô�'�����TuCx�|}�L�����'ZŒ�v�o�ݢ\�����A�ƾSA�9O<~���7�t@iOU�{��
�+�1��P;���N:�W"��2��nOK���3>���G�]W�w�#�_�u{ޯ�Ԓ���uBØ�/ k�x�ɗ���oPGT���޹�"u�
{Wk�y:�枌a�uZ���7���dl��m�u�����KB�oy��?Q�ӳ�z������@��<�c����}�8
�#�^jɁ���#-�)P����017EM�Ć�Uh�b�gk$}����xf���H��5��G{/�����O90���.��"hҙ�v	X��k��_ ��FA����U�6�@Ի;�_a���n5;���5[9�qbwsV���ب#�Z#�z8�my����ݹw�"u1�U¦?jе�{w]���w�^�y{bv'ޞ�)0�����|t]׫�eN��䛻�d�5'��U^��M�w�1I��Q��_�J�΅1ݛ���:&<ku3�[�X��e�w-�ߌ�﫵']�ǲI�����'��~N�o�!��A�4�����w��Վ�;�Ϊ���8^jd�p�D`����i4̅P�Ow�z<������=0P�kh��N!���0�z#����ۊ*�����sއӽ�zo�7Vq�Mb���qY�%���tg4[���{6MJ�h�;[|�됓�Q������"���s�}~zw�"1p��Q���B#��i\kR@X�p�ۼy�]����`�]q��F<���2{[�9Q�?=nx��F�z���"m�v�܌��=�{6��G�{+ζ���N�����Ok�@��&��O�NL8��7�o�/:�b,o�ʜۥ���:h�}��Y��l��Z�sL�i��Zw;?�����@~�@E �������"x�����A��w�)Ý�9��^��#<m���\��v���e��lP�^v����5�Ǌ���p�x]����3��%u֖:�ҬT	��	P6#��M].�����Ek�Zٱv����8�8�jW�52�#�-n��8d����W�l���ČG&�mq��ky5t1f�*Q�-L�nSI��TuH��n/�1��h��)QSE\���M6f�	�q�b���]B�����t�n��Q�.���k7evڦ�p �.�6�� 冡MP�..��b�6��E,\ᘖ�Ͱ�%�(�1�6d�vsqf�-�f���4H:�a�Zj�m��X`3�蝻3R�f�F��$�ZȶC��ki��u�[k��UEqvRRK2�5��Itڤe�I��f#{Z��L�إ�iF2��Xԕ����6��6�v�9�4����ey1��w"�����1�I�eх�B��j���)6��wl�D����s�n�tlZ3DR�s.s�7��*X���5�M�ImEwd�ah
gmU^���s.���<iM�J���7L�eA�%��`˝M�jhM� ��bj1:�HG鿲����r.ޚ5��!\�M�bU�N��b[�n����xA�s�=�<�β{*���d���>~�F�E~��*0` �ڑ�����ڈ��ivs���-�mK�V��z�5QS�ˈ���1���'��M�P� �����|#{��gP��0�9"�A�F��ń�pI T ��Cm�*�%���2�a.P����R�H,��pwG\i��}�y������ړG&@f�>��
3xҁ\@P�����]���r���d> |F#.�(�MgsQ?iAV�cw�	�d�78�.���B�6B3Q̇(	$�H�YUR�
[�o[�^;��6�,Or�G�OP���.�i�)���م e���*+r����a�4b�P�ˉ�c�&v����4�@��f)XAY��K��,�׋n�(
�qYay.`��6�5ب]u+��#CJ�M6�e�7��9��$/9
��k �(��� �*,�-�eAeH�
�Z�"��<���Ƙ71�m��ƸБD0Za4�&���QWέ}�c��*G�Iխc��3�7����Q��}��I�Kwsp|#^� ��K�����v8�s�X ��@�֋����=����g��I��ύ^�S�flҳ!K$��tr��B�X��"u9���� I����Va曄T����p�vu�|��T��F�qx��Ң�6�k����6��':��Q<Ƞ�#$YY*@DJ�`�����%ds��9��OЏ�\8n	S����0�K����P�be�����Or�#ᘄG4�ɆbL���D�����n�}�̜
 ��m��6Twt"5�2�Bb@�P�Ord�Ow腬3s�ۖ��%���D,6�s��Q�%���
3�ݡ�qm�J ��N���� �"���m/���}#b4��D)RD�6G� H��zg%�ڣd �M�EZ�"����Rd�X�����;�g9{�|7j%�]��Nj�F�c�#";l숂ShI�a���q��V0�}Z���(!QiT5M ��MGM��l�K���*z���=�7X�B�|�
$ZϾsP;����?�Jⅸm#3�"��B�o�6��0�lN|4��'
zݥ� ^�Id�ng�8���:���m���9����4��Yv�{�PU���$X)�`�E5+��~���m�����+���'u3�?1v5���Xi��q+�]E���\J�_^���J�{�&=��j$���Q����L�)㯢]��L82of�� �9
U�rk��������E6x�� sR;|�
(�8ր%ق{�'���)r��}uR4M�҂��I�xO�ʮ�o��'~��L����N,�Y�@�E|�@�-����3qe�ʰ�Cb��pZ�X�22휷Vm�t|�����*��1���S+��e���lZ��l4��*�h�L��
�#�f�Ħ�6���[�`�X;3P�L3+��m���N*LV"����-��;�{j˼�qܔ�tt�&��B5,���AT�8}x}���O��Ր��0K�(<��B8TkgJ���獶�8d�&��gN5 a�i^P4�QfP�-s.3�|/b�\0��>u�Q���F!"\��߾��[�������Ol����c+D���0��e]�� 鵢Y�x�B�o�� IQ�j�����2Ol�v�2��t�H܎�qZ�#��3)����g;������o�?|HP�	�T�Y���7���x�����D���>,���P:m(e���Ř��� j�\/���e�$����B�����נ�޿9�u�����g,�ε�]qFWD+L�&�%�@��Fkj�0-[�	�������>��af%�c2��f�#Fp1
 �+1����Rt���\�S�0���S�� ��
��ͺ�T���j��V�Sf�\���6�7��2 ��'�R�@U �PP��,A@I:e�É}�a& (H�|� 39�m�O��D��\�nP��+@q�\���>���2g3.��cv�%k��Q
SLs��d���[�a�]k�Q�J���bd�Y���c)��q�n�H�P��O.�V�WK<T����tA,M�c�m�0�⛜2�f���[�$�ǝ.�@�UM�t/����S��".3�((�x��
��hJ�ŀ��A�5A6xs:ˀ�޷� ������Ӝ���A���h3jm9��K6E�Mh"�W:݂V]��9�Gg�9�;��2S.j��KciNc�D�t����m�5�M�����4�?gp�S�|j��ǭg�~�O!���eC,����%�ҰɊ莫�2ɳT�Y����p�o#;�D��9=[]n�^o\*���f'���t�'Ah�I_��R�ͺi2�[Dhf�63t�#f�nMF���i�s�6"$�R�], \�gJ�:�X͊��+��mW�ė�\�:��Q]6�r�4���݈c:���5a��4�W4
�[������K	$/-���݃|��� �Z��Q�AK�ǳ�[б)�[�W׳�!��>��Q"�R�"�o� f���;k�t�p!���Qk�%�yO�8\�@h��^la�B9`�5=���A@�O��^��u[.����}�O_�sl��	�:���Y�����9˥1�ߴ�/��_|�a���,��(�Ӎ�ˊ�)W�<V���cc�<y0����v�$�L�u��S.q
�R��QoW�l��	X",-��,��pί�w�S���p�ߡB�bL��b�з�#N5UG��P���D���q�J�8ː�	bN�Dp���f)f��o��=����Os赾AኸM7+[��0b���Rf����p�|>�w�Y���

%��a��+���Q���F���ofn�>���z,�nP�74��{�e�9��t.bf��ژ���ﯺo-���1tQܱ�5$d91�-)��}6w�VR��a4�1+q\^�f�+XP�Ѭ�N�X�uS?��1���ص�sz�c�UӞ45\Ҡ�c��d=�S�Nvó�����T@�DKfjn�3!�q7mC���"��g���$}�-A�q����Rg���M_)(ĭƷvi��.Ѧi��HxO�e���Ǉh�{$t�w��\�!�M��'�DeQ*.�����tP%����ݢ�J,�t:���������z6y��|�dv^�{�<�O���'V%��z���+1f)��I<��Mo0���EQ��Hsׁ,V�y7kr^[�s6�T�v�Uc���ѓ����:�����o#�"{w�Y`�ŲT')�Y�6L(���J�<,���K��f/Ao�]���CpS�dB%K����B�:_�5F���[�5k`L�PR�ͷ-߆�7s B��[��˶n�Rt�?^Xf�,��Tio`*̫B������
����)���(Y%{���$�>݁.� ��s®����X�^�I�~�񥢍X�����bE�N���Ȗ<�Z�ǩ����4�J*�CHD��0�c �4�TQv�Xf0\<���]�Ȧ_o�4i���>b�t�y����~��Oe��pt�{*Z!�w/}�e�niZ�=�$n���,��{���xw���-̣�m���H�LNh��9p �9�󼇯���.{���^"�@��� ���p�B��
(�,G� �TM@���:�e�m �VM_İ�g�
��:��@�
v�&��q�E���;��ɼ\�.�1�Mί�3�dA�N9�n��� �*_���I�/}�־a�����ge�sMFQ4w���:v�xv�Haf Vo4�5��~�̛'�N��G)����k�K���'H����C�C�b_ԕ����������8y�ո��T뾬s��sf#s�b�s���*=_[���=��3��o	Y��X�S���,�
���'����\��<���c�9��]ݰ,�b���2��ߚ���K斸�*ߴ�~�@�a+�1>9��q'~b�=���L�=�&�V��~C	���i�+~�2���~��\71چ��w(m�:����i����N�;��UNO�+<�LYS���s����d8��4ɨ=�ό�73F��2�C�J�I�����+7�a:�`q����~ܺ]�8Β~�M}N w��ÐϷ�n��T�VK�ۊ�b�Y�Q�N���幃�\u�K�u�69�a�@N�Fc�o���kNN�+>Ͽ]���� ��E�Iϩ��g�Md��r��[�x�����ݬǪpTL�\��[�D��Pj�Q)�t�ʛ�`]
V�s��EQ���6�8`n5���X�Нe2�]��ݚ,K��e���Y�����r�ffi6ЛU���4���R�%��,���W��q�ε&��J��-��!Ma��j��h�h7.
�䏔,(�u��ԒX�Rm����e�5���suД�1�?��aM�]�n��V}���q�I��q�5�ujE*��aIs:7s���eA�{C���f�E5Ŗ������C�a�{�g�n����@����)�s�aw��
��B�g�K�l��.䫪���� )��[7��֬�H 혛��SQ �T}�����
�qU隶����ߛ؆P?0a4�P�uS3Z;Vݳ=N�ω��g3����,���rv�5����+���p�Q��kŁc8֪��9�N�Z��ؕSXdeܾ̣\u�]@��i�����b]7qy�w.�< Q�[J�j�Zʗ�+3��5'�Rc5'}��I���~7��~�ܮa�ЁY�}��8��m"�!!�:��f�u�95����K�j�%ِ56�Un�1��vb5 �zd�$g����8ʗ��ۭռ]ddu���q� ��n[�G]�k*{׸N0=!�_��j\�r�X'	�j�J�+��t��s�y̆K2K�*�q�v[�5���es�e��@��Ru���@������4�UL��Tx��� 
j8��ݮc�:O��3<�L����~�ό��6� 隟e"�I���{�κ��Ǿ�>����f4����am�T��-��֌��N�l!Xy�"k�%}R������h�?HI��ɨu���~���7.ݼ'���2@��:f {�5����5<�$��(c�9��yM�w��:g��W�		q���j�ݎc�=�%���6��8�ĿEt�M�BB�R��,���A�;���w����;�S�n����9���tv�B�W1�]_s�񹻗��,֫}�& ���:�p��fcpx�n ��c�j�隗=���f]�:I���j3�&���B��x�E���w�69�`���w�b�*Kɨ������[�G���~Dy�#������^/�*�Bn|��B�2
���Ϋ�P�"�`���矽�^��~C�e���"Ϥ�����@���3��t�Yߚ`�6�GP{�و��`�
���~z����b]Z�6�k���ݕ���M/��'!���K�"� ��1>��%f���k5����F9�\u��sg{��tUdsA�}�_�	P<�M@��>��eN���P�b:�:���.d�u ��-���`��B�cWG\wc�I��f ~<�WnW0��'� �{�}� �j��n8����qk��~O�?*ڂn�	��R��̩��K� :u�Wp">ŵOT����e��5ݡ�ʈ+vk���nL�J�=e�g1"fb��F�l`$��$!�P��!�Q��E�V�����+�Mk��i��bm��Llն_�n�i	����tK�3�\��R�M�&�ԳX۩�k]2� 8s���r	[ƣa2G��됰sF,p��{�!R�ŕ�t^L΁��ܩ�֜����	��d�m�����<O�9��gW�)��ח5���L>����Þ7nc�>�<*u�.��ɨ�|�_�cHg���8ʗ�p��g_�� 5���_��i��N�=�$$9�6Ԋ�`�\�T�un"���Fqx.�YCb�J��hb��uݸ�r�Ĥ^9�jHq�y*���V+(jU�J�t�)�:m����u�8�%��&3RzC�=�-縘��dlelv�^%�\���S�wo36�;öt��|��
�u����:�p�Q5A�f#qk\��xI�`6'�? ��~� lH6�w�A�r����U�����{�N��N����:9����)����?E���X�qz��Wܷ�H"\z�������:eg�~�q�I��f?������-G����5
�u9��w��R㮙�P�tf9���Xb-G:�k�p�E��G19�����bbKɨT���%��S�:�Q�z�q�w�!��}MCY?����f��ȣ�u��������:N��w�f.9�'l��{�YY�^a8�0깳��-".�����n"�\y��#]̴���:eK��C�@5�Iߴ�q �����Ӯ2X��7l�r^�u���F��qY������xXvш��6{\�7PpB��̈ɘǱGp_U�}��$��"����"��������8ʗ�0��H���9��״)�{�98�^'|L�cQ�\G�`���fcp�<��;srt�Y�}��e~�2��u͍�03;�1����ØG�;���(z��xh�p�sr��)6C#��'''f���-Y�'�����ɬԞw�k*]i���XBqY�{��8�8������qs[�Vt�ߩ�Ђ`�y�s ����oT�X�f9��N�o]Y+&�P��@��<����!'lԹIY�:�MC�:���x0^*���Њ�ǝ�5���d�5'��e`����w�Ê���	��j��&�'��c6~��]���QU�6%�D����������5���w�z�ni�/ �<ϰ����bX�u�@�>���g]�k*x���o^��0��ۦ��-��Ck�&ڢ����x��a E��*�D/?b�@ }��S�z.W�`7
��܏yT�?_� fЉ2~d{�!f8������X�v�i@lWE~�����y��� N$��q���}���
ϻ>�n\�\9��;�")�^��x�و�Z�n ��{��t2����񙛼%]A�1{�nj���P
��1��K�Ә>�J�����x�z׆�.ne��y�����7���P(�뎴Qʣ73±r�XY�m
������^�T����h��y6gn�\HdU�b�H`q�H�Hx��pT�8m�؉�q;uf�>��|��`٭�1��8e��fNk����)��9�����^���VN�nv��)����W�q��+���;l�����+��o�WLGr��;u0�Mȹ���yj��*U��T7
(9B>�T�Bt���n���L݉�ݜYD�Q�M�e���ی�?�M{�xJ)����z�F��F�JfSN"=$�c�
ВȋiS�h̝��X:׿n����jW���l3�t�ݕ#|ɭE�t\ޯ����#n���Ҙ�j+�A=�v�D=w���=�	5�����x,��k,�
�{F�noFEI�2�*�]\Ȧ�݂��2���׎
�E��� �_��}�Q��X��Պٝųv�m�ȶ]ֻ�l�`�/D�hߴ6���JZ�t�6���vhm���(o6�e�Ť��c�#w�@��I��`�``ul�S�X�nɱR9nWR7] :i�[4�`�J�t�e Z�t�=����ɖk���7*�]��]m��b,	)�|Ue6]�MCP�����.�h]�-�̥р�T�9��:�9V��]n�5�(�3(8x�UbT�Bż��-���T��]Ʋ���,�U�U[)�.,3���2�	���Li�[,[(�t�HZ��3B4�ز��f`kc�Bٸ+G��4Z,��4�U-���ݝ鳌�	�<V�&0h��٣Y���%�q(L��`[�e��1���*Qk�u��:��X�s&�f�鞭���e5kE�Į�D��]���iv��&6oQ*i��7�K�u%Mj�00��D%��
06L���j��4<�_:����T4�]��.�H*��5�tp��f�	�]�G&�rn]�)6�cu�Xͷ���f�6�%��X9l�j�鵙[�cZ谥�h�n��k�*���YY���e�s�]iW�yVy���&+��P��l](3O]����ݗFyM}S�Z^.��W���C1';�����a�ث+�;�o_��'n<��"�6Dt�R�dFqgYIl>F���{�� ���G��,����	���Lӣ'�%�LT���ulx%�{�����x�ue�1��ӱe�ϧ��3�������+��;9���X��y�s�'ޓ؎C�؉��Û����,����H@jv�����T���OLx��gy^2F�t��cwX;ʑ�֠�7���^P���}�Qk�R	�Ǜ��^P{ӱ�v��X�.f��v>�i�s�A��Ē���F�ݥOu��{&�����d��6ɼ��fc3Bk"2k��z���/��Jb˯�2��%�3&�H��2g	!0]2��H����Y���*��!�#�.����B�Ϊl�M]Y����!sz�m�KTf[u���KPlgz$2;u����0�XkU�ʱf6���	I��<x���Q��.�3Z[�2ܗ,?N��s|��Tu�OGRI���Q��ⰆcP����MP(���w���@��O�:eF���g~i���� ��{d�jN�fʁδɩ�Q.7�o��uE��@�j��j8��h�q6�E5�{�u ���a��7g��u&W1�	�تo�٨�\`�
�w��3�R��;��ԏ���s�3��ߓg+���~p��z�����]�L����Tw��4�-�E�:`���ˡ� @�����K��S*��ȁ}]��:�GQ���s`pu�*�8[-� Y��C�o�A��>�W��罷�\�����&!�\���q;���ѵ{5��q���T��BVT��a��af Vu�wt��m	'lԾ��s������IY�O~��P9��;8��Y,kߝf޽�v�������y:eC�r4���[�G��5�3�ݍG�'��q��ןk�i��y:@����5��Le�:�ɬ�N�1�y�rI)ޤ�}����=��&�[[����ѵ&�(�}󜃴�̰� 6C;�+�`A uzD�w�=@韷peK�ߛ~ܻ�)5�$��s��tZ&`�E��q���cP�?a<����?g~z陷q���~/� ~�����LP��[~�lQ�c��8��ɘY�5B3��S:�E�*�P�)F'4�\�n�hTili�Y �H-b�~�����>gĝZc*Mg:=�;�\��N�w�����8ʞg�aq�;��JL����:���U�n�rAO�X��u�����[�P+<�=�S�I��^�}m�h�Kqv�'f��f]�X�w���������=���d��}rq����$�1�{I��=w�n]tί^Dh~��n���СWF�� $��65���Y绁�f!�xx��>S�qx��-G�;�uF.ꋻ���ċp�;���'��Z�un"�\w�������i�̬�Tt�כR��;�,ÝFs�p��t�
FsB�?"$A'ՙ�rMeO��|\���s	�t�� }R��\2q��~��eN��%f��?{N������4nf���wl���T���h��g�H�_4����d�
�u�MeO�P���*b�k1�;=�滅Ó�
�����N���~�VjN�i��ϭ�� E/�}B�gܻ��5���q�LC`$:�N Vy�{t2��X��ӆ�����|�o�����M���b��8R%Ý��8���'�k�m��1�tɨ�o����#1�?A��� ��!S4����3��#�&Y���#�(�}�=��s��F�-l:�\;�;��m1h�(��YaZ�i����6�G%Wk
�074�5!b��M�X f�3��[4�v�׼l�È7.�騻q��Xe4��Gf�l��lW;fP��tvl�	r�s�v�!�46��;��LJS�	  I�z7�,�ն�ʢ�Ps�mntr5���ӹF��f3|�+;��k*y�Y����C��Q #�v~
Npj@~Dc���<���t����j：�u�a;�@;f&g�x�����&��\s��w���ޙ���~�>�אXn�G� h�듌�g}�����Mf��v��w�c*�ߍ����N�+>��]���g����$��k5��S�q�$�o_g�!�����u�����JZ���-�R[<|m�,7�:gl���&�Rui���u# c<�=�S��_q�����O>��@�Y����[���Wv����,�����h��325��z��
.⓪�qI��E�VTY*F�}"�|�ɨ���YS����%�����Ϸ.�s&�P7��Q����"j$�`u���uvw��5��A%g�P1�Ny���z��CT$�RGpw����]ހ�$�v7`�u�1���9������t�f.�f����P��R1s-ë�8�i���H}|�-�{�H 
�?��#V�g/���>��>�ǟ�0�6�ֲ4볽Y�Zf���zm��D��b��$��Z���f���ze�kI�R8	? jH�v�1]�w�N�
�M�wZ�E{q���C���I�U��נ��r3�^��<o�+��w�����ʌ��@�У����k-�-p]�I;@3��7�T]��
?k�3"w��/���;� ��vk���6#����nNo|���/��Ԣ�e,����������8+u>��~�P\��9��k0c-]�Վ��gq͉�C�3��_m�{��]$�$|(�>DA@PY�^u��u��ᙷM�����}4����>ͻ`P(k������P̰�4<�-;�n���w��g�����g�v�ӈ&����H7���oN Ev$y�iē�nm��"
i����}����Qv~F�2gܙ���t8C�_�Al�����/�u���{����!謎4��8���H>����	eAp.�rsפ-�g�_=*�/b���H�V�!�n�M�3-��r6�5I�L�9Q���L� ��h&�0�ki]�ܤ�V���j5li
��f�9WT�)l`-M
�J���5o���A@�qe�&k���˝�Gf~�r��yrdl˲k��i�c:eu�9��%�fD&�m�v2g�~���]F�a�Y�\�-L �����wɽ!�7�`Ƃ��V���4  \6m,F��0�`���L�&iW�#~���zTá�BS���b�gGI������ʤ ��%�� хƤa�]K�l���#����e��z~�5��+5�<���^aҚ����y7�q��ƭ=G5�iJޫV�F>�BA������Wdt֌"�*0�d�$����7Z�W[�
�4��7`����
���"!VD_�/��pްڎ�
npj�0�� #gСgDD�"3��\��sp���LÚX�߁��7"ay��ʵ�P�� >���0�~9b��ڦ�FW Բ���s�>y��JjlW~DB���_����� .���f�	����R��)��>�t(W舟D`G���ۂ�q�T����m�FM�����
��&,3u7dO�/*�1�o�X�����$�}����5��%-�u���U5�Tؒb�Z݊5Զj:��B3؇��'I)����x���M�k�w�Ma��|P~�>ӾZ�,��晁��ІPŶ��.D�k�"��WM_OJCFn8<�N��:~��pO�\�&�����uL띪���|!q%��.������[n�k]yY\�g�S'eX���U�D%�2&q �]�z�����ny^���
cr2���ԉ�ڪȡ�	;t7"��'f{.{L��S�Oz��.[�
4ɻ�w��m�>�@��`�*Q��h�ί�۞��竞�F;�vk;�"7;	qR#�\�+�{���Kz9�Oyِ
,`룙5����6	"��Ь�_{�$Z>\�u_yh�֦:�7��)�\���fj�c��׾qh�~
)���g��և�'�)�Ȩ��g�;�τ�5��c^���b@Gz�1�<�/e�tC�lo5]��Wt��c׃�K����ܲS��0�,�U�t�'�ә!���R�X��"SZӓ!;��������L�Ps�n����9����#3H�F{m�����<~�I��~���"6M+����I����K��G���#��x�P�]�]�.��"?r��	`��(8M[Q�z_C���YK1��sN8�k&&A9	�m�Z���U嘖�$Q(��֍9�^�kZ�ѩy5/�}ڹM\�9��?��B��� d>���up�#.d��J�n��!��x|숅o5L���3���_�����Ӟm�V*��}�����Ƚ��V�����Þ�r�Z�
xDG|.<���bUH�pkfҖ78,[�m�$w�x�i�A6�č��7�QL��	vtM�UK�����Y�~��5/��KZǆ����ije�G�  >��X�
�,Ye`l�ր<�«�s/�降<i�f���sy�#g�E�Z�t���so�޴���I�q�\�u\f^�"H������W/*XG�a0зo��S+���q�J�DB��o��'^�4/�
@2��)fG]� -��V�޹��Svۚ�M�o�L�A���>�����Q�Z�̅ çK=��f�D7r&V��}���_�[�\E�F��D+y�w�@_
���
�".�Q~%w? fЈU{"eZe�Ȁ��0��B.MU#����/faW�B������͖�Z����\c�Ӟ��SNVnۧ7G}�r]�/J��τ�ov�Ͻ.��������9}�����8�bl+m5{;���0Q��[������tl��,�Ye��]b�xf�:��񱌉�h�j�W1��V�4��1��i5b:��[2��aLX��6�֮tҩU+1�$���-�^����	�1 ̇������7�N�����=�qP"�y~|���8X�Z`���W�>>wbDB��fU"�S��qam�`8$��kϼ�Q��� ��~��^Q�vTӈ�*�|����F�qP"/���S+����C����o�i,�S
�@|����o'=�~_���a��CA-�Q��&���v�ܙ�+W�!c�S(ߣ��%�DGf
p�A%T� B�\v{ի�qu�ۖ#�u`���Q�Bb�vR9kET�z�	���:o}� �~���dJ�ˊ�����Bh�ڪG}dF��jDw!��6�u5{��؅Օ�!O�uUW�g��>�4�jk^yLK_�*}~�T�2�﮴�X��(���A!�.ڬa���vu+{I��v�bOx����Q��
�?>��U��O �����^�H���+L��^� S7�[A���÷K}
qDp������C~& ^L<y��ۮ�q��vѓ�b���[Eìы��?�?~��BY���[��i��,�7`�+�F�4|�UN`>��jJ�n@�]����b�Z�Q7!H�{9�
 ��m��v2�!�tahi\V�V:! ��՘[�p�6fUyo�L��׻[D;�E,O�~sYB!s�)�oѣ��)��u�v@1SK<�5�șDǯ�&U�]U�������*�iv˕��y�jv�����Z�"B��ind؈W�kTjˋo���>�G�G����n�ӆK�B��az�#V��W��f`��+����+*+��&bX��a��̫���p��3���<B!b�'aCF��#��K��S(�a«�ߠ�*��O�3�R�Y�#e�ȉ�}.���2�~=_B�CmUX�5�
�fe_�F��ˑ0���[iКV��\��9�����P�7+$_���gr�F9�T��]:.p��Ӻ�5[��fE����ϳ�֍\�*131��V6�i��B��,h���E���e��V5�Gux4��̗Z[�m�5&Ef�Kim�:\%f�I\�@Â1A�T��m	j�m+6�^%j�]�:fo�$���yl�!
@�)ں��͉L��
�q��������6>���)�C�k���R��S���P�=3*��@�]q�3���V���¤� #�"ak�S(�,m3�C��w���|��Ȍ��n��>Ҫ��� 2�UR���^t���a�F2;�&\7k#�Ze6U3�E2#�q �bpل��l����2�G�e˸
���pj�b�^�ާ��n�3~��E����^��U����;���X^���	�H4�ffW�Du=��Y�bKa���ibe�@�Ͼ���Q�C�k��2A1S[�����W�"�F}���U�m|`8$��\��e{�?|�����̪�����lpE(�@l�IEf��as��K�6�,]�l�I���闯yL�ǥ/n"�������(�Y!.���]-�CO��{�D+y�cZ�5�d�������5AIY�M�j,�\��9��a�{-��@����B#��� |L,���â���)Uw��ޱp�"!Re�uȘ���\D(D6���ҡ)�ة��S
�B��������E,���E5��g��c��͛Z�wP">����~�x�
��c(kIT��(��Y"f_�"�_��0�hU.}�2�l.��.��2��!OAK8e�U��}�&]�b=r&=��q�;�Y����l�X���WOh����z�%FubU+�OT�����H�#�|Qkҍb�i��Bt�f�����qL��-��V���߳��y3h��[1H5����\�56�aR��Bջ�@�V���~|��&�O���£z�}�+�裒à�g
q8�'5q��A�b�/[��V�S35c�<���.�����a�LL����>�������ק�/�Z1V;#n�T��z䵮nm�O�����iͽ���UUdz�믂[��Vk��<]Zt�p�ό�j���o>7��dϦ����9l��7=��k��]��`�Yqt��򸳳�d�7��|���@՚��=���/rƅvdFh^�_�.c��}Q$>�W�&M�u�x���;j�mq]Y�&;���mn9��Ss[
����݋횃O����F�e>���5�=���'��<�!x��
i���W7ͫ��"���*��UgZw�˩��H�]�>��ƽ���/�	A��i��=��e�A��s���
[�Փ�������Wxrݯo��^jx��o�[�~z�'>�v��5,[�����^�}�XG@Nh���V��P�ۚm4@�ڳ�:.�;�N��(7�Y�a�t4x�`K��+���k���qC(�ԇ��t�^^"�'`׊|�S����i}@8�	��J7bd�nUؤ�3	�s�V5�gD��l��S����%B(�GX���55���my�(���R��Z;��b��R��mJ`�6eA�4h+[tÐ���L��:��e��i1��e��)�J��2�Į-\B\�Z���c%���6f"41��I�]ͳ[c4ItA����!0�U�Z/./[K�"4`�R�2Ү��16RkTk�9֮�ae�b
�v�t��c��6V�bG,����2kXeml5a���ol��#��J%�k,��aY�@awX��:9�Ej�˃-�*i����LCXI�oh��ck��!a�chR;Tؕ:�maV2���,2�sq,ȅ�`hR����R;�6`��t�ѵ`�f[K#f�-+Mk�����aZ�Mc-`hi.z�Bl��5"T32�+�\[�����ńJ0�ړL����sG���,B؏8�*ٞ4YmѦ�,TB��f�^�ꈤf#3Ը�l��DaL7UV����حp�J��Tpcl1�`F�lfj�6ݗfqYA]r�m��-L˗*����_���>���'i	�{#.���m��z��LCCl+��{�g�Wxx��y\ե��[!����ѡ�g_��Е'�z���M	��C�y7=����/a�X��0�/,����26e HE�o���y4�AC�q-Ы�D`�;O�'G�Xw���lX�P"�v:w�C�m��u��8{w<1��h��)Ʉ�CZ�,�c`���Y�[rC}����	�����.�w��i�}�u�az�rl)o��
���w����I�ry��oB�����#��ڦ8eɽӖ/6�)���{��C��=
��jX)B��ݢ�pL����1�Et�٤d�-�uvkKOc˼r�����LGB���8���_t.R����M��.u���j��D�<f��]כ��2��+i���)�bcLؗ4b�lc��:������ȗ8�*Y��������X�m���+�(�A�Ĺc��6]ti���[� t	pN�#�86
��mpHXm2�BCg#f��P)+�pMbs[�>��ؙ��Bi�%�?����PX(E�9����Y�x>����"��A�O@�$EeGSs:�7�B�e,���M�8&�<꽙���Y��hʬca!�ˈ��K���yx�o~2�Xķi�Іѕܰ��y�t fH����.���Է�!M�ϐ��N+
���8��,����
.���!�����h�o�^[6%;��&�}�	���Ka�;nf}���8�ei)�ؙ�c>����۲�S3����"�y�7��tF��PgI����ؓ�߻���\��y��?���g�(pT`��p\hX^n��=���Rd]�[ޙ������S�
���!�F�`G %��s*�yE�E��;t3a�8%����F�̘����U���R�d)��i�_f�TױΠt>�����.���vp�+��M�@��R}��:�̺�����[uW�;��^l�S�(�@	?Ee
�}|��j"����ߑ�.DJ]�s(ߡ��Y�V�M��`�b�-M����`[�g)Gib��ͯj�Sp"�8 �bӕ^Go� �IwzxPΆj�}K�P�|n.��٩{��=p�)���a/q/��7�mz��t�h�8ܨ����\E
�7�ۡj6��S���[`��.�VĢ��7|���y����
(,�A@F��
�B(M�����(��G�{`D/���5L�«�߾d$����V�Z]�0�L$9���8���ꧯG��l{��<>s��p"��x�P�mU#��iQ�S2��!M��/P��n�*:��������*7�r�ܱ5��U}�w���`A�n�dP��r&���P}�³�M�/��:�W���I��O���We{����5��^K�ݱU:�g��&��_]�ۍ0�V9��\-��(�7v�)�k�h�-^`5���h���b�v�����K�R��&u��:8��mFZ��F��#,5�e�#f��\�p�x�M�&4��Q��B�A�ڍl�L�3!�H��`#!�u�����\��ywBgD�	eδU��0�3 �[j��e�o���W�R�Ps8���q�,�{�G�;�X�=O4�.�-�!���}k-E��~�o:"�ǖ��d�����&dD*^����"b]��L�p5T�z- ^mU/b�;�M�r|���>��c�2�,�-��n@D��j��]Wߞ���(ˁ��׀i眘X�Y(l�b���G#��s�ʈ���ʎܬK�+��fh�v��yي)f�ъDYwL�7�~@Y"����~����k����^W����S*����y�S+ؙ��-�%�o�{�2�艶 ��*o����M�<>d=�&��}tA�g��l@ �$��0��)e+�96+��\�r��x7�3��3~O�������>
D7ڞ[�� 	�كw艶0
"]{����T�F]���Y�]f�湋�&��/�Unk;[�k:밉+�/.P�ȻP�'M��Zb�U>ºfP�W���}�#�))E��v��y{/�r�u���<}*+ ���S: �@�D�V�刡�%SKآ�\����̪L��f��Y��$�Q�i(���x3�ً���z���}�;���\U�~���Q
�JY�[i�����瞧�\���yN�)��V��q٥��[j#���Ș]�3*�1��`�F��"ec�S*סEs�펱�$�7z�R�=?9܄F7�<�s�n�̪�r��u	��AZ�o9�[�^�n�@!�,H��>���ӣTX��};/�|�\"���{W��MlY	���؄ �Vl��(Uy3+ֻ�U܁�Vr:ḇsj��r">�F�>�x��C`�&*i{TB����g�eZv��q����U���Oy\���
�fg@d�S*�g:�*���2��Èf�B]��U���z#�n)z`�''_�y%��s�VV�8��og���Y���Z�;{���m�ɻ뤒-!}i��A�n6�!0��e�e�TL��ܤ��E]v6,x�ʡwRPأ1��Y������7q� �i,�e��"�Z�73Rҍ�������f�$��4�fڸ�jgBU�¦N��ӂI�I9-�ν@ư�(�)l�jp4.��	���h�Wg������������3	��̪ލ`���`ټ��}-��G=_N���t�+�Cj�c�uns��Y!/u�=	Ci�U�淥¼ٙ^��x�"\709Zƚnf�&^���2���U3�
F��h���5�WB��6�+Kf+Y����J��=����lu�}��U�x3�mBa�T����7Ef͈x�Z�¿']w��;N2-,6��f�	{X����CW��>  �I rEǜ.활{�`|6��N�l�-�*���2�3�}r&��2�q+~D8-Ӯ���誕آ���A����ˊ�>Z�]�"eH��G=_L��d����Hf� ��n=t&[��5�FU�\�Cף�����K>�M��T=�
A�pA�uH磇�%�l̯b�R�ϸ�&�ȭ��M[�����~�"Bа��e�����bԴX���K����1��~<��k�Co4ϼƙ�$إs�����u�=sqV��O�=���~tu���B�w8g{��~� ��z�;˵5��v)�d�4��.I���Ws(��r.���m�����+�VW�"������Q�gR�=>�)�Q}���ï����>�(?a<w�u�*���~ʆ���JO�����䇌>��-���w�kN{�/<qN�(��	�7�����o���U@F���b�}u�Y�e^��r+����<'����{s�f۽����z��w,WӚM�⧳N�P�Z�E�چ�>b<n�7a�;¨x��]��my�P��d �q�yF�#�{ө�<#�	?6���=�wm�����S���2���c�o�u��n���X��4X�WFo�Ym��{H���c��-o���5QG��j�)h�l$�� Ʉ����֩Z�d=���V�`Ť^8���`��+sN�r��C�Į��o�ܪn�z�N��������3v� �#hj�W��6����/�c�[�z�����i�{qU���B�+*���k�xN��j�����ʤ�[D��v�E��ny��=��y�p���.yJ�>��k�����hƆ��P؛R�#a�U:ed6�CŃ.n�POI�}d�ąi]t�Gpnn�zX�=�҂�n���	Q��6rS�q�;�����&.ͦ?���^v��hYe�ɤ\Scw_�=�C��j�tSº�L��H�:`�ʼ6��ڬ���,;aJ0���n"0n�y������@l���oK��/����"�() �������ͽ���|a8&M{��L�a������;p]�c4 �	��������,�r�=3+֢�O��놭�v�fH�Ѡ����0J8pnb�{�=T�2��P-n�W����.�,�O��O�D,�������a���`Ѭ�,�s��g=.�L��/B�mUp���"anl�S��@/x����E>�9.|F�[�ft�����"K�]8vJt2lb"%j��"H�"9��$�,��\pd��UH�C������U/b�]p"1�|���i�4Q,�w�C6!LM�4�q��nS"/��>�w�dB[�`	�o�´-k-�4�i{w�Nd}��4� ^���P�hU%�Q�C�>�~��֢��JY�[-��?w��be�@���o9H�KIK�!�u���綦W����jzJK�y�e�j��be���sټB�V&�X����C����T6�Ճqf�ޣm�($���@A�V"�fԊ��l�՛;�`pжi��-6�(�KT�� �2ٙ�s��+��ue�B5�X��*EM�n͙Z��U���0\+�c�t�L��+pd\݄]+�u��,�Wnۘ��
5�-pR���,,���B�B%�%�>́�Z�U���}��n�M?l�=��r�V&\T���C��h11��D*��߾��aV@��lo���;�������3� ]3.GL'�m[�(�?Y"e{=3*ף\��d������a��^t^�z��,
ij��F"�b����̬�S~�4�wkڢ`�tnb�{}6�-�Y#�1��a/��44���k�����x�kx���\䧪��k6Q�V 5;��{��/W�����@k�[
�ս�UJ�Q���k����[�l� X4k�g�B"Fb�[��?}��[�s��f���U\�5���v��\jøX4�� ـm�Da�X��f\�T�Jm]��D*����]��e��*��ƚn��������V�42�\�cZJ��yD)a��%K�^бw�.ɯR�P9D��G�h53��OO�{���X�Aa �.o�s��e�
l�4*��c�U+:"W������evH�:e
���̯}�-��>�2�|�F>�^f$Bb-��fF�0ttB�m�qm�n��{�2�TB���2��fU�(hd�Z�Z�ﾳ0��L��D)��
���	6�J�o@�WY3�}XY�c��D�#�jl}��C�ȃ>N��@�������=�"��(���F��$b�Ặ^n,\�ibFП���KeD�^B��I�X�*ł��!��N�o{�!��<�Ǉ� DC�z�J�DBφ�^��+����l��X�2�k��K,I��(�'�(�W!~W���uV�9Y��hA�0��^բU�~�l̯Z�~�T^VL!2�ޙ�X���ӓ.�b�W��Al*��{�UJ�Q
�F�gUJ��a���a*5���de�����ٓ2��c���!q��h�Ӧ�2��Α��׺�fs��GAkxʼ܀l����lJ;Am�\�s+��ff���qmɄ+�i���#6#��m�j�vW��*��c��(���+�3�7@˰iB�E���,�ͨq�3SU�RX-r�]m�f5���Һ�*��H�	'-��ʻ��u�6sa�#�˥`�qs��ò�|�W�/&k�O�J�Jk�>�[jO���Y��숛a��{/�oRM��s�:KG��Ԥ��e	KCb�+&��H����}^�߾U�E�]��m�y{T}�dA�dG{"7�3�*�$� �B>I�R�E3t�3Zb�1M��LQ�� �0�~�>��֠߼Q^<.�=��֪9DTf�їw,���Qb���L|��69W�a��܇�ͽ��}��,� ��X�(	��	���ss�3���������K*�smS�YD}O�1;fg��Bm��U]��*V�ʯ81��Э�"C��i��6w�1���"��ab�Vn��;.�V�T�\�%Vh`���E���ɕ��Ir�� ��ͫFQN{�0 ��^Hg����<���p�P�Uy{����*gN�9����{a[)9l��gn�U��f�}���T��7}R��A#�A��dX,c}��n��w{���]ͣ�8/�2`ְ���q#�������27�� �Ț��\~����M�����F��еim0B����UCe�ł�MELv����?�=���γ�7��<�@܍"�ή��+��C-75�b��=���o�o*�:�3�����8uL��N,|^x��ꊉ���cF<�����;��g5+�����|�w����AV"�TQV~|yïٙ�{V��מ U���3�q/�; ���Rnkc�L��y�Nè�ו�������m	��� ����8��t�s�^>��u�l�ݨυ��H��D�n�����a~��f�񱁖��nhg���/w#)g�x��}x�l��7~|�����R���C��v(D\��֋��3�0��-m�ٍ���P�R�O�܌�CF˨��q�8�Ҏ���B��Y�jqa!��1�C�����蓼��8
K0�Æ%�;Q�%]FD�j)�c��l܉�JF
o\�	�T�ü��K��7ŗ�����t[�E�œ��-� �fX���,��XZO���m��J�sޗ��,+3v5��ví�Vd�{��wk���t'n1�Xvb�`��k"4��p�^���oe�wtf*X�e���u��l���Ș�,����e��)����t��tq޹�_����~�B"�p�G/�"'����s�J���{�/�����ŀ��X#��t[�;'v5�1�숸�3Vnz`l���-{��ڹ�o�w�+��|���k��kL��_��ɼ���Ũ���`N�$lQ��1Fu���=���COZƪ���gB]ItnΌ�Nm�V9��Q�^��Ls�"�p7i��]�06�Y@2n��i�Fb��M��͚k��E�������d�hm5ecj�і�s@�4B7Z�8���jU \��[[� �M�d.�\�ti)s �[\`n�\SWCp�6���:���47V[4K�q�a4�ZV�F�驱��D���@2F����#*�)-E���k���е����JP������C=�Uo^M2���;P��t�R[�vL^IFX[�P%�u�5݋4����M�Vaౡ0\�-�Sak���ƀ�,�D�JL�]
�`5��Ƃq17%̺3Z�&�R3K1�;3���4.��7�1�w\�ڰ�eb�lZFg!3p���G��C��MMBƚk��v��AR$��:-H!s-ڑL����0�[UU��V�#�[s2���L���&]43�u!�F���7"����lp$@�,�6�II��s
�8M,si���X@��g.�˦�K�#X욡rgfw樬L�9��l3�H�M4���)�2� (525T�NK��p�1�`�\Od,q���fԡ#�n��pH�Z�&�Ȯ��U�݉su���S�7uC��sQ5�E�6��K�&�BJ��4f�%����6�PU�.x�Z\�7J9�A�'+���#��坧]|�c�mN��='^ʆՕ(\������0M�99; �:�0挧;v�/`�F3q���Y�h�<
�bզ<Їe��" =_l��U ?C��t��>���Q�A^Ic8֣�-	W��}1WP_�=w��7DY����x�kՏ�y{�����]�{ݨ5��oG��u�j΀����C�s�FX;��>>��Ɔ �%F/MbJ���/��eL$m6R	��KX� �tN�21�ej�v��T`�������-��ɹw4��]����,���N�@��k;5n��y�z�����m�5NT�bk�ƹݩb,m("�Q̤�n�a�Yd�nk&���]0�7q��j�	Y`�I��VZ�eKCAp��:v��hͮ�-ؚ����$x�K��G1�L����q�H@$ڽ���U�z���]s�Q6!�i\V�1X&ulݨM�ͿC�����C�����J{�K>��FQO��L=�������j��*�kl������}W�����r��'}��ޠ<~=��z]�����7���tb����JgJ���M��3j ���z6�#��?��g�85�`�_�,g-�b�T,����ĖG]i;�",�E;��Q���VOo�_�����gJ�,��"�A#����>��&��Ϝ&��U��99��~��^.�8�?��Ҝ v1���Do��}�ŷ�(M���S�.d��?z���O�_V{u����cWA�w.��U�܊�Jo>����Zc޸��S���^���L�����ڌ���W���c�R6�(A6[K��2�l)�8��7e�W�1܌�@��&^��ӓ��A��4r#�2���< ��!��R�m-Q*:��{��XQB�\'Q\ D}ޑO9D,�c当񱈆<1��o~�Z��l�\F}��:x�	�(Q�h%\�l��ap#�v�r��U�{�g2�.�Qv�
�&!�@�'��B�ȉ�zg-�c����ш�GW��oG��hD�a8�� ���B;�"Y�ё�ܥ�5�=5{뗘,��֋��N�d*�'*un���{:%w�=��;RV�U,b%��e�	 �	��˾,d&U������ȿ�^��K�՟[S�.V�˩�#����m��st"�\�G{�A���o��TY�����5G�������sM�ہ�}*���ł����Qy����w:"k��S0�5]�ݱw A���w5�D=�Z2{�@�ک��[<E���~���-"k�e\�Q�9��f�]8���\���\fm���*�[�!�v�1�0W,-͹��l��6�.���Ĵ��.�;J//0f�ы�y��y�j:�%��7vXX�Jh��B�&��B;Fm��s-��%[Nԫ3��G�+�SC[,�4�λ�@C�jJ ���[amV4j������}oL�)��DŚ�#6�uZ�s��/��k��6`�I��P��Gm� TO���}9p�w�D�^��Q��,��꼴�[q�����ĉ��&�s� ��0miuM��k�T�����\'T{}��ٙˈ;�o�*�qf
*'	|���r�C[���=����l��y��B=p��>��1d�y���u[����'R[v������Y<�'�����[<������g��.�s����_s޿_4b'�R�RڌkQTJ��Gy�k��κ�	�{�zb�J2}��������b�3#|U�[�Ͼ\�\]�yQu��n��ta��
���#���=�<�^|
83��PNq�.B�X,��!BQ�s��� `Eߖ�r�=^��L��w���a�O{c�	V����H.����k�_�&��=���ȍ-m�M��S�~�hS���'"��S��Ѳ:����񀓘�#㯪Ҵ*TZ�-��X�+D[�Y��ϻ�y��r��b�Fx}���>��|^�U�D�Uix��Q�꛿�����L6�)Ay�5��q��݈�:���h���n�#��𙤏��6�R�<�=��m/*,��^Tt�8�Q=�������d���I�o�C!�o�y郶���Dx�&�d�޼%�Uw��܊t�FO���mKF�^�rL3�W;qU�rk�w��}[F�TT��QU��i�v�a�-�<��L�zb�6�0��z��&��[+�D�vC6�l��w�1e�^���F��vY����!�kF��0�9���c�ϭ����7d����u]�3w��}*׈smȜ�3
�
S���c/'��3��"MX����/���)̟Jgi�]A߻���^��uǠA�͛�xe�ի���& '��x��YW�`[���z�%N0YnI��b�����HU"�f��l1���ռ�
�^�3B���3s��L3i�P3y��B��jl���n�r[̦*d�j�K5��K.ԛc%�l!�vڪ;U�mm��w��m�JZu%�R�X��(K�Ѡ�a��1m��&a�,f�:)KG��X�̈�a��G��U�}c�hT}���;��������Α�ğw�:>Ll��N?"�Fp}����R��$��z�β�O�,������CmT�}s��-��R��R�2�F�f��K��\��U*8����ׯ��ڈ)}���$�]���۾��K�Z�b��.���$E3��O%y�S�y��|��������eH-	A�1�өCG�����ƒ*���Y�RK�-�i���K�y����@�A�B��7������"��{��^�������B���qr�M��4�U�ߟ^�U��d����Ir�Ap�n��"�]��grO�H�V
dV!P�|d[W�n�X�\��K�O'��so��9J��mvy����P3� wӰZ ��1$·�Ff�%M��mN��d=Ѳ��w��79C�̡�z��t�N橩
�	T[������\r���;Mb�~o�^��t���i��j��K߁��J�.�����0��h��xd$�tf���dU��,��RV(o<�N�vL�=7Lb	�ޑZ�=���:\�9�g{�}A�����sd{u��=t#[~B�/t�.{�ȉ�nO'��+��?S7���V�'~"��th�V��Nɍ�2�1*H�ߠ�
�f���Ɂ5�e0E����^L�ٰ����b��aR�Ov�z�.�k�g�n����w��E�i��q<�
{�5��$�y=(���͹AZ��y�+M��e	ʴ�1�^��9��E�X<&#@"�I��=��y"�Ap"!�wd��	�(+v瞊p]���� 61���L9�囱��K#��R�qI�^�h��E�L2m:�ka0t聁����l���.FN;Sn��9��ۛs�#�wM�ɦᕬ/*:�;��O9h�F��S>�{�_�8��i��[�5�iw`�}+[r�J�����Ɩ!�:fQe�Q]Y�	�ܼ:޹!�3�֍�H��q�¹�xy�Dgq+�:�k�Y����1���c���B��@~�q�k�%�-�2���u�x�'<�}�l���v��xf�a�,��ꚷ	�6w[9�s�N����{�Z3��wFȷ�F�yR�b~��E�V�O��+K���qF8B23��y2<�Doou�<@��X��Ek��&g̂]봡��'AH�:��_<��~=P�֥��"*,O����V��+�ߋ�RN|,�]c��c�2o����A$:�uq[Υ}`��>��\�7jlT��M,�j��T�ٶ�̦1�����f�zw�R�������}������ك�{c�h#�a9K������f��F�K�������ȼ��:�r�Ǎ�M~�3����=���u��#�w�3�x���y��}�Kh��J�PH�A #9l\���-�g���ob�w�����~���@#a�Y,��r�j��M��ڵ]��=�������[��S0�(�Z �U��*�������)�ff ;z.��Sړx�EM|(��6�G;.��f�*;���us�Ƿk+��ʑ�Q�[�hL�c��,���x��oR��)co����z����hP�P�$Lp�]��,4nZ-f΂��t�k0�)��m�4��YKт��%�8��ne���M�&5�ҷL��r˳�%���&�8�D�jb�B� @��j�A�\�efPu�͍}8�j,�V�XJ�]:�סsCov�%�&�d�!h�r�pf��M9�ğLx5]3%��-�;y����������EsK~.wk�Z�/��c��
6�|c��$��]Lm�{�P�*wq��� �ɳW�<����R���Snɜml�53vXқML�"՗c8e��}��}�M���gV�P�M��l��2&6��D�Q�?#�=���{UKsT�s*�a=3R��$>�O�-���Xa*T��~�?=W�ߪ�*g;��
 �tx�P�6��vt	=0��nǅ�hr�����@���1�o��^���J�PDU6�Ixt#wj�.�3�["�����Lp����V�2��͂��v8���ɴ�����S�w��*����v�[�=U3c,U��v�7�8�3x��R���mXm�Sވ���j'螭���"�RB���^ |��QU��?B��-h�\F{���p ��oa"�
8�_��w�lͧ�'����Bߨ�4��	��FKkp�K���ɵk�H��Ͼ��a��\� q���_Y�w��UWc}�
�=^��z4	�ԉ�$�%�'��2���G��6�5Ԓ��'�~�2��Q��L8�ѯuFŘ��ۮhn{VD^
ӡ���YJ]Øˮ�u�F`�d'H� �@�1{N����n�a��ٙۑdlS�����A/���"�[utl��\��K��Q�[n�<�a�^�5�fDf�Z�	$����j��7��9l8n����3a����#~��e#����`�L忝��@u/pn����iV߶��n ��#}�[ֳ;�y�}�=�c��j��%�Df@��s��]t%=��j&�MZ�ܣ[��e�X�8�A�%��Wp%��U�!<I �����	����#�r�t�YIX�m��35�	6i6M.&��)�EeXX�WF�y���=�j�i�\�Qq�]���>d�� ����9��jS4��̺j�!�U�nmv�q�X��a�V^U{���fl_?"��v��L��F[�1��
i�i�|�(Ϸb2���&r�"sܽ�(���}:��Gy�ex�����N�'�{
Rm#�}us;�{�|�߿_���.R隵��M"J�]6L�bl�m!)�z:�^UDz�f]�g�K,3��;�S�l�d�>/:�g�&b36�f4���X� �^�-Q�k�r�L��t�C���3��?|��a�Y�|��`Y�d��-!�Z k��ވ���-���>�ma~�����eȓ~����8u��� ~�蜶�a�5�0ω��0+���i�F�.`�u�h�eP�5�oR�*'�!�����|2�uW�=�K4�_ME� Va�MC��JN$jj;�}�:��`v62J�6<a`ۤuNi���*k�]�۵}x�l�S�8�ayv�?|>~�K�"��5C�N5A� ,|b�̟Zv>�[mQ߮�D���3��Md�>?+q�_|�>{��ҭ�h�v+��k\�mt SKPel�h¨}}53)�{�&{�}�� ��X�����,R���;)�υ��-�v �{�3}��bsp�>���AFpyn�2��_��ש^L+�����֤�pf�?�H�Fz��߂b9���^����p���>G�|�����^������a�#�g�fM/2ٯ��aY�a�����%�8�Ƽ��0�1��q
J��jj#}���������Q��M��(2���~L�͠S��D�B���^/�W�h�h�{TH��"�ozg;J:�#�ğy��&0��y-�1;�b&6�;��C����W=G!�dF���4Ȋ)�9{�7ݤ��g�y�|�+����uwl�O� ����[NC�7-wK1�p��t������{�����	J{��' h�+ޝ�W�9�c��7��R�[^�ϼl�ǰC������{C�\�\����,���j~����m�r�4�E@F9���)	��HN�ɳ�����4�l{��P@s��Z��g/+[���nW�1[8����p\s%>��Y�z�no��[|�i��M[�X:��B5�WULo*����U�#w<��Ά�������?i����|�MQ����N���8un
Z&�b�o$Ğ��뾝��uۨYF�Lj��nUE�*�����1^���D�v�w�6�F!��@��GV����@���/I�_Q�7�T���w�w(��>�������9��M�fI�����D�9�V�����J�4���!B�i��������ڈ!6��smb���kn�ML�]��SS3$���Iv��;CXSDmoh�nlB^�	1�iF������L���%�XUk�ٰn��5F4tc&ntV5�k�lf��v�Q�t!M�%l�n����gWC0U�;D��Wu�B�+V5깲�]JEDCYs ��]IC�[�k�f�*�)�J��h2��XF��ګ-aV%�34t��e W,e�`��B#�,36��4Dv�#�c0��(�f�[Ns�Zx͇U�*h�ͭjXvZ\ڸ˥��Z<T"1�ه&��#�7,XƄ�ufk���f&�5�.�o	���L�º�Mvf���8�c�uf���<�-&�Q�vl��Vi�ڑ��F�:-�]F0�r!�� ���yhKX3����������&	H�Ņ#�96Ⱥ�4�,fNԳA+��5��YYL9\�ƃ���a��4)�ƪR�p�a��u��f��M

:Q�-*��+.�mZ7M`T&��R�Q�с�f2�h���fj��+H��k�K��3���3�U�J��W�r� gg�W���g���?���i��nA�k̻���6M	���>%�P��]�0Row!��x��[Y�)���֔{�9����kЀ�k�"��D!�����7�����f}1��pa�H�Ԝ�Qn!�m�?\+e-�M@d�e]0��yB&)���,�)����0��/�7�p��kQ�r�߀|3��{p��=�)�<�I������}�qC�v�ӛ��{EA���=�L����K�˕/*�gm�l(hTS*��P���X�2��NS���:�d��k��P�P� f���K���a�θQ����9�#���>���VB��*K�ͩ:2�!|�id� ��оߘ�)�[��O +l�DA�gb�sh�/\���n��G��n�"�� ��t�vf�{�D�����8wA�US���NE�s���
 #
�n-���E�s�09���;VԏY��G��sGeB�jDVbˋ�Xpne���� ]
h�.����2՘����@�C0ִ��eX�h8ʨ�[ي�;+䚬�	aR,^\^�͢��˳�c�2:-c������*����6���sd����8m��x,�̤nr����R����i�g0��߀�+��tEQ�-C��KG�-���z#~���'Z��^/��&O�3)��n7�%C���h�0ei^�K+nj<����o?"+g����*W�FV��a�b��S��T��tWy�l����{Gc�1���fBQ�*��jb���,�1'qH��@�������M�4:p����G�l³�5�;i��|σp�V����?L^�D� �f=��c
l�肌��#G�mA��N�]Z�_y���JQ�]*X뛑�t��P3F�9NC0Y[��l������>�L=�0Rs~
�g�����5Y��4��>��]��Z�pe�� �����p٫+�]S}A��B;���=�~P�y@/������q{���m<k��8��`�y�v��X��������������>�}� �	��CI�&���&�+kc��T�&��ZbO���q��#-	�k��B���"^?z�g����Y��2!�l��R{�
�9M�A�Z:
��uZ �@��م���ebrfL_l��M�ŏM���!p��wV]:��u�&�U�u��R1 P�3~{�����sm-UKZ,}��Fw�g��a�^��n""jf�J�5^���4��M���y���"k.d��}� B��>��\Nw�~s 3�6c�����kpr0�UjfV��n��'}�˄C!'G�ކk�7 -��VX\σp�=���Vk��0��L�iL�F�^睺���ECk�s؀�/�3sq".�_�{x6&zf���2�H��-M@��1J��ZسH�+�2��̬@�ىRڬ͋��u�4�@H4)�SBm����K���*�a! �����e��
���Ŭpp�ЩJ7h�D�іEֲ�ts���e��w{�x)i
pHJIN�<y.��]��np�6�B&-*���:��73K߾�B�Lҟ�j���������� ��A��㝁z�0� �IIč�C�}�Lv0������V���\�t�J �4b��d3h���8|3 A��0�]�~z�~������Ɓ�&��U��Q�ĥv_~���ޅ�����}����҆ZbO��\�.��/Hg�,�`��^6�F��{�t�;!�EN�a۝�t�;w��P"��
E�h�qx�KgҞ}�Y��E��n�"7��H�=� �"��Y�8m����D�̥@u=@�Z<ʆ�w~���sfM/� ����1	�D AeC�k]T"�fŋ����J�cf���q �,b!]o�Z�8�G� �u�^���>��� �bo�b.�s���M���.�!YW���r/�l���Y1��ƭ�h��7oa3��<��>Ak���ZR���wL\_���FA�5�|��Sg�;���3[�L�		7�DHƙ�7K�E)`�b�؈�S�BE�V͝b��#���2� n�sq��c��>�}mY�����3^|>����l�_���c~d@IU{�fo#F�;^.��U(g�	)�d��n;��ܩy�r�c�0�~��E��t�=�E�8�(9�N2�yۢ�݁���P�R�k�;�x�m �Q���;}I����D|Ǟ�����!LLe�WVSr詅\�\$V�b.�g���K��(��X5G؟}����Y�y��}�(�|Q,����y������S�
'��|7b2�R ;ZƑ|�Y�8m���3��r#Y��׌&G��w,L{���3Eŉ����B6����ɏ�w�痼�,��k]5��gd�ĺ#e���<��&4��`��\����$C33`q-�uvQ�V�c��[�kYn�s)+)j�\M����6 e�\��GYfX\�%k����X�a��5������E��*��*��*��:�H>OF��(�P�X�2����L�:E��L�(=�k�� S�SC<8nI
�t���!|Vp8�8g����zP�C�������ȏ���/�?�x9Q+o�K1�5�G���y��~g���1�طj���H�X*k�[*�[>��6�g�����XY��x79�Ϣ8��cˡH���9���n�Tvf#����ѱ�7Y�k-�ms���?@)|>G�~���U/�g����=zz>RG���Ix���K3m�[g�D�V�����2�^ �A��Lt2�FM���}��qo�s���	�Xa$!���m�#��諕���ʶP�K0��q��I��3\�q���Ă��<Y ��ܙ�bp��`�!���v�Z�)�菡\&-�\b��}J�����Y0������.,1.lә�5���Lm�H�p�p�̸��)�"G�i�N<W.����7G%7ϖx|�G��h�w�=7 A��Eo=^۔g*b�w=�j���<�l�@��\<��{�>�e��Hr��S� ;47��}O�1���ɉ��=V����չQ9��-X#+R����r6"�f���qlgRݷ�����⼿
�o]��݋Fޮ����2�R:�z��=�
�=��v���h����Y��gh���͛����7wї�vN��]ia%�࠳F��`�DD!M=��(n�
��6�5<-�4��ڱn�"2�)�g��=ʳ#�5��I@�.�QY�&S|���O�w�-�:�guȷ$��{���=�h3������[ڨ��w4�LVm��;w#7	�fr����X��<�P�� DhEB��JX�>���Y.��A���?"h���:zn�j��F�"���xt$g5��L��������'�N�mt��n��� �II��,��<x$��n���sǖ,=��G��v��d���Ϧ�8N6�DȔ\��I�p�e�K��떙��m�",Uc����0�\��'P�%��eED��|*�b���1e�#eF���(��d���*`�4ᝌ�Cd+�U��o�:Q��	9��D�e�Gz������ٺHW�@B�����l�Wj�	�ȣAi��ܻ�G�]�8����۞R%�eɻ!��#Xo�i:DKEf+v�iBq�,d�e�No������ ��?{w��}/W��]�.�/؜+1�O�b�q�|�@�������;����gI:����m+�na��]k7U���a
�ъ�ճ(����Fq���v�Ag��0�s�kw��S2�\s�)��%DB�Y�W�2w���߲�9�j�<���WW��������}s��Ks����r�MՃ�u^�ڈ۝�ۘ0��s�}7x��Q{��k�9��8�u/}V��H��\R�"�B�o�۫�G�빼�|ߤ��4�͙^.��>�`�!��E���p�0�-�WmuFh��W祙��=x���Dm��(�QBO���ҭis��Iw�[B�����D]lE�����U	���;��TY��E�d:��>����3��ʣ�آ��ȣ9����tbn�h���³6����ͽ�M�Nr���f�tf�p���룜�A�R��p[�M�)C�IL�h���ڐL$l�9�U��g6�@�,6�ۨ�Ri���sPn�$��s�L�l!\&�(Y���y ��.��llf҆�89��V�m�n�d��W�Z�.�9nc�P'��HTU �A`��z�Cַ�[����n]�^�1Wm���m��ԧ�z������y��A3|�^������s�>Z���k��r��"��s�Ǡ|}�b��h�Iv {v&����
�q����%�����]lW�L���h�C��!�hD6�	l] Д����(�9�stn:�b����#��+������
S~ʤ���ި�-��sU1��WzS�Y��p6ʣr9s��p�2����q	�����a+"�Ш1�AaYD����׸w��3x'���"fs�{��|(�yW(��䓁��>��;����wE�����EypȬ�븚�/�| Vi)��lY�Ŕ%�:+Zk��	�tq[������3��8C1'ُG̉��ا���'o�8AD2�g1gѭW��E��)����;�y���iq:��.t	TN�tE�_�y����>(���+"�J��(����`
��T"1T��U5�ꌡx�\2\���*�~�x>��B�5�D7���ڹ~c�hDY������������3WRaU�.Xdu�������^��|��y�m�r2�lI~� 2��ُ����x�i$�_�^3��|�&����ȇ�:>�ػ��c��|mv{�����u��,��un��`�z5S���r挮���O��I*E++������XQ`��޳3<�Jz��ﬁW�;WT�}�|� �(Q���:�]E���fX��	Da��{�b0��/����c��G_�˧��ݏ@�x�CG~Q�7r������n$��1B��t9�O���3�|�q���D�=ɞʈ�a��Nd{e�M&m9�纠�x���dF�\�	번=Iu�%�OOK��<Ԭlx<��d�U�d�ʷ�;+[�.L��ˡPc�%�s��5�&�r�7�٥���S	[&���9#��ti�X�ԃ�m�Tl���V�cm��*�4��-�;c��E�`�J�B��T���6���R)*� ��AJ°PX���(�������^�r�WW��,c��gW2�.���~Sz�6�<�rc�lA7�%j�"{r;�9�/{f	�|��!��^ZY������e�mX�(�BBw��O͋�u�p�.��יp�wG�7�|7.g��=�+~�+��ϓ4�*\�׉�łʥ[� ���D@&��ڒ�O�~H+q��bg�!�m�?٧3K�w��%��8�U��wă�P���\�'�f,���Z\o�gUdvܣHͯ��$��$��-��)Z�!QJ�PJ�ciF�kB��Ұ����B�����/�y�޳=
M�d�y�-��G����һ�sECJYdU��^*1�).�
kf%y�D=H(�v�o�o$I����|9'�S}�'ct��B۴�����i
	qn6��r���_�ʘ��>�Dv\F����ğy� !*9�R]�����b ����o.�/mL�Xߡ�J����˪H���K�D�3�_Z���ī���Ȯ�jhu���;�,A�,5-i*�V)QAIQJ�D*V���U���EdZªV�B��Pm
�dY*T[id������b���-�!Dg�،T])�LO��h�D��3��	��^Z�l��,F���0&Vc\�\#X��"⚅����k������3|�;����p
'� N-�S��_�J7��B�;툫a��z'�N����������>�ȘR�����E�ȳ�������~��jU�v��A����7O9��H�N޿D�	V)@F
�QPD�E T��XT+�FՀ�%HVB��3}��Ù���$�6|>�7��5��{1#�B�e(��h�`3gi�-yp��jp�wg��eDW��K\ٔ:�^
3^z�E�������"ﱳ��&UV��o�g�O7Rr���fs���q^�8���I���%@i%F��WN�y�{���x�~����>$�#I�I$�I(�P}�(�}�_<_ӿ���-�f �e�Z~�:�3.*(� �����!" 2"�  2*"�� "
���*� "2(�f�UB@IT�AXATY d@� P�Q8�%���"()"����(�"��Ȩ
e�
��C j(�R�(H��D!BDA�fZ!�(H�fARE	 ej)�XZ�AB
(E�d�@���P�@�Q��T !QD�U��A��@.�"!pU,�\T	�@��@y�~����:�X��1�!=QI$DXA��Ex������a�=~�Q�����^���z?�?������ ��!�:�`������:0t�C�����Q�A��?~>{i=^������C�'�������>����_�O����؈"�m@E �_�X���c�������p�څ����/o�?�u�'�S��b(���g�D�0��ȴ��>�?c�T>Ӏ����
(�s�U%g:�:�!�>>��h�1��.��|:��@�$D��F�B(�`)(��X
@�$R�X
@��BH�E"�(�`)�$ �$V(�X�A�D�D�A�EB) #��A �$DH�A�$E`)�DB(�P��Db� H"@B(���Eb�"��$H
A��DA"��$X"E�$A�ED���A�$�DF��$Q`1 ��1@��Q�� "��@H�A
@H�EH�@(�F��$Ab� �`	F(A`	�@"�
D(�V(�T�$Q"�H
@F(���E"�X
DF"�P � �`�`@  � H�T�$PR�
AA`)A��A �P�D�$PH
@��H�ED�A ���Pb�X
AB(EH"@H�@
EH�$P�$(�`)(�"�(�`�H� ��$ �F(��$ )"D�$b�� )
E��b�(�X ����AH�D�HD�H�P�HD�H$ ŀ0#*@�@��"� ��@�H�� A� ���DAcb 1�  ��1� �1$A�A$@!0`0A"
DA�A�A"A�`��A0A�1�((Da"�B
@Rȡ ,Q)�A � �$H�Ab�H�b�"�"�"�"�"��B*���$H�@"�A!��`�XF*"� ��AX�AB��$D +ř��K�����m�8g���p��(4�@B_�zO��=!��8|C�F=����|���?dt9�����$�����ϙ@,�A�~`��}?F����0����m�?8}D,ON͈|'���a���&��u$�z=���=��<���@E ��(�I����:'����o\���}g���UTR�x�����F/�e�'�n/��!����>��to�<�}���ȤA9=A�HA�x� ��)�y���#�-�V��e(��+ ������A�A�\<���O]�DP`���?�P�����>��w��L{y�}49�/��>����Q=���?s�sj(؏�0��{��� "�zG !������fϯá�'a��r�$a��Š%%��gOs��h�����^��N|�.|LmN��r "�h�;�*��G��x�|��9l���C�""f߻ͱ�g��r�����y�("�~ѡ�@��? �2�yy��P@=g�������\�쾈�K��񼆃����_���<_�rE8P�&��