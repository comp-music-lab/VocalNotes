BZh91AY&SY*\��;W߀py����������`���            8�( �U(
��PTU ��(@ @ ((   w�
 �)���{���]k9���Ӧ�m�y����G ��C�a��pW �ClQ�ktc�{��+����ouP��xuz�e�-�S�s�h�ѱ�g�m^ػg����m�w�׆�і��a���ɭK�]%J� 
�à�z�4�.��9����g\��6��SN�	
 ��5�<<����L�f��u�N�4і�Q � ����n7l���2�q��:d�ݺ��4�G�ڊ�^K5�MtkBt�N�4靇���T���7^:k���:��a��z� ۣ{	�)�4::�4�]��            jy *�j��(����@S��jR�SLF� �# CL�eRM2��& G�b  �CT���MUT�        JzH&*� �`&�dd�h�� �4OALMG�����S'��W�����y{yv=�M?$��$�x�=T��B�9%�����G7��]M�C�bP��O���q��>�t���u���8�U	�q��_��{7��^޵J��=�^������L�20nm��;\���{��6��? !� �G��H.>�"O���o��`cV��wDFɸ4�X�4K�=�SI�w���Qv�0��������b�֍^ ;�B�XŘ�1 �4��5$���Z�����S;Q�{}wG'(J��ئ)�P�˔фls���5��ڷ�75���8{�:MTvN�U���+��W5��j�N�� �kf��#�7)���0Qq���GXѝUޢl�^����ԉܸ�
v�}u�)rk]#Z�"�R��}�)�K�zb����7#շ�����B�׿"�8��&��WYgeY��εG�ou�.Qn��z/g���.C0��x&�#s5-}�:���W��:p�=*���n-+\d6L]xR��s���té��B�6���:n�L�u`L�ŭ�
�*��й�)��4e�
8���9�n��k	��xӺ+�"�u㨼��i#n)e�$��f�]��]d���Af��7����wXŎv�ք n�d)��;�9w��B< |���Wz637�����[��r�ʆE=��L�uʆ�Y"�+1n"s��.�D!��8��
�ʰ<��I�;=��؊�� �{S|:�rv��1�ڇ	 8HE{srk�dNπ���B)	��6T���z=��Ȁ��Nty3w:?�7"��v	�DX�5g�٠��'7��K�Y��鎞�ǜ�wA�mzX�Kt����2m�n)sC�/r�k�{,��ww"1������b�������2d��Y;d'6ϖvxn��V��k{!ާL����|K��G�bO k+&�ó���L)�d�����9��ۆ�Q��pM	�#ܨl��ݽ�o�*�'J�9]wj��Gخ����x��4�n	�}~�N��S�(��eۋ[[h�Lq�Y��m����n%�./xRՏ{w�U�:��݆�]�n�ٯy뽍���]7&�ส=��Ln�o+z�8�G9-����Wzf�sr��vfr=2�7�`B��Rm�n����׉�� k"��Q<�r��7��^s�E�q���Ӂr���Δ�����A\NÚӱחD͸.s�z��⻻!Ôb�����7o9�� .���·��gb�Ʈ���wI���@�ɜ��ΗK�	�cH������b/ZF=͝g"e=���;��-%�ۣ[=��p�o�Cp����祠�Hn@�5��\���hN�sL�[f�|a��%wi%�(�:8�qrp��w�:wo&P�0os�5�׷��gq�"�����V�yI<��G%��]+����1��d�΂�``���M�(��5�=Û�;���n+��oE��1UtM��|���1�[	p��zX'f唕y�ʖ���7��t� �OD�gnq�N,�4���$#����O�s9��'y�M`�;�ry�lݘ��/lm�Aj�d,4v��[��T����ө:���g������XʹL	���N�;ȳAǿn�NQ�`���'�rؓ���ORn'I�N��$��E��"�xA��Aî�
�����B���@�C�5psK�ۚ �.���ɝ:u�&��}���t��.�-�h����0�F�sO	���N��v�<	�7^�Tٳ/qZeܱ��|���W��){����h9w���J��s��Uտ1�4�Y�����+ćmgpYY��e�A���V�=>L�٫���@��A�쯋�]�����5���8���=�H���[��s��s.�[�V����UG3ngg�v2��������͙���G�ݏ,��3̀2wAɎZ���Orgk�r��y�d�[��`�b4����b�6�Cp��(U+UC;��y*Vph���XsA�)� $�qb&�I|�۫(<ogF@�����ǋpgu��sۓ^ș,�dc���w�E�!�9�l�6����+�ba�� q廒i����vrFt��u� Pqh��p]�F��ၐ.���8���d���Wf�;���]�|.i�gV�� [x��&���Ri�V�'�yf�T��2�Ov�p���`��L��kr������<ĸ�¥�sj������N.h9K��	�G�1�fIr�h���`{��Ǜ�A� �o�}���<W�N��h�������Lȴ��Ɨ-܄�Q�20ZU�uɌ�����v�U�Eȳ�9AK��+%�)��j�ӂ,���R�3[�y���t��m��ZW.sl�v�5�҄���K�9N���!A'��9�>	��Z�� =�����5;;";]��J�N���U5��ܾ��w/�9�� sK,W����7N��]��`K�I{R��i	L�m���7�������~A�o���ly���D�~��!B�����#�\�li	2vJ2�]k3���.�q-	F�,�/R��3�0���[la���	t1�� �4�2� �֚�:���f�=a��&dhc6%�����.�fkؓbЙ��L�i�P�m��8c�v�A�P�Y��34%t,%��b!tAq���*��&Т8QX�f_+ϓkO%�%kD��feqX�ۭ�k֎�08�SCGD�ihY6���R�m4Wk.��͆�b��� �K�h�#�`�m��ͭx��)��Ce��K�Mn�Ɔ�J�U� JU�����y|[��yfZL���G=EL�4�4s��qk���f�[[��Wl�-�р�̐�JZM�w�����ڔ�,�b�*��EΈZ�S[��X��l�fM2b�U-m�����h$;hJBJ��6ɤݥpc���|�<��sq,�
�KlQ���q�[a��SMQ�p�3�YV�K�V�i��VP�Qe7��V�ƺ�* ڑ����kc�Z٣�C%�n�	X�hܔ�����%�:f�J�e���.cq��W6ܦ�
F�Dc�6$õ�y�e��v���]�M���-l��Hu��ZE�[�r�LF�Kb:]1*\�И���n/09�2��&a]y����U�4-KG;8��:r�+F�[%�e��h���I�.Ԉ�M(��.AՉR�;9
1���INv	N,8�9)�1�F�E�u�+G3&f���v�ckċB�\kn�RZR0;Rn)Suq�&�Ggl�Z���c&Uv�t`L�ƶ��l��!F��Y�5�m�٦SL\=s��ti�-�����E6Yh\�m,3hŮ�٬Ϋ\
Qư[E9���	�s�5n5�0�P��j����1ZQ��n6մ&sJ�f%���K\LJ�1�F���R�j�b�u���@�%.�ʕ,o��k,e�^Yw.�ǰ`��o\Xn��L����f�W����˵{3H��(]�,��)Ֆ��(4������8%�ΰ��6Z�l�V5��r��Tt�-��C��j���v�`<a�u,%�l4�ƚ]j�6Y��^&F2�C�V���-�շ8t�a�ue�.Q4j�LYNk����׍n���D5;6�+uw]p۲F�ˀl���Y���k*��6ް4��ɴ��<�V��r�pj�*�vr�f��i)c-F��9��W�P��i���m"��\��h'�������+�hi�0��{[�Դ�`�\��yX�G��ʶ_�`kIc�����n�i��KfŃ�X�mZ�+i+��R�lJ�v��K��XIe��U��n��n�7F�Ǝ.�]rJ$p<60��Ml¥0���#2��,�pv,�.׌F�`Z�`�P ;uKz�uUt�کQ��u��q�&,ri��F^���n��F4��7R�<>^���+,�;7TCCP5��[����t�)�%ӉJ���T�ոx�u�A�!{hK^�eg�;�a�Зc]�0\�(aJѶ`&�ֈs�֙���Dt���&*5�4m@[t�6�3j�oi]�fe����Z͵ێ��k�����X+����2l6��e�o9��al`ǖc\�`�����R)]�R�S-�a ��r��lQ%4
�i��Q!v"���!\�J�uD.sa��:���WJ�]L��(�vѡ�eka�g�7�6�	KsI�c�a�iu�U6�l��.�vɑ�n��)����חR����s����C,b��F3]�a����Y	��i'I�N�{qϒT$�:�މ"��o�����=����߷�S���T\���S�(�K<]��^���0��ۏ<��o+�z!|}�c1��F+�MPBr�&M�&H4�jץ�r�g�������	�G��ܰvpR�͑sUԑ���������P�-�,X!x"��Đ�z��gsYq���E��c�V7�TV���!��y7��-{>���v�א����˾���3G���gy"7$f�<�U�^Z��s6�ݔѰ׵�`Mѻ6ח4v�T��o�}W�P3���G����v�7�.:>ʯ8k�c�B��8��{�Ǖ.%<���˾��վT@u�6�x�y��� L�ѹG�メw����c����>��f�4��z��^��U��a�r�'@��f^�)��Ȭ�ype�&���}P��fX�qL^�J�)���	rԁig{�5�q���I��s�����j���uck}�H�ǻǹ���άv���ô��޾�1M�V���z��	0�J�ב���=��a>���;�.�-�y�<���i&Q�Y�k�\���ݧ���zv��т&�ݛqh�����p��fKP�	��D/y38f�O��ᗷv���|�y?|�9���iq��{8�9P�F�{�G�� Jq�B�U��3�<�<+<�@�Ư4�T`\��k� ��j�q����yW+x�����FL�74���}�@����Q4b���s�+���1���^	23�!�5�B�U�5�F�9�w6k���wG$���o�٦͝�K�4�|Ϣ�}=S�fg,��V���������{�}�4����)��-�<q~龳�O�W�9��eٹ�S==�g�nE㫷�T,��y�:�i�&�޻���dOf���c�d�D6[�NC�V4��ڮ�\�}�=�]���m��8O�su�K�EkW柶.����;��q}p����m�f�di�������xI��6�{8tO���F��%�' ko��uy�GeS��4'�M�S��}�뤷xi��o�F/p[�������ﰾޓԲ��<��o�;+z�j���������ٝ���i�����7�^Q;Fُ<�,�tP9�ӵ�to��z,޸v��4�s��S,��O8iZ�7�&$�_x�!�0�8}�&u��{(�C���� ��Sٞ�ob�E{e�K��/d���q9�(�^%7��ҳG�mQqt�=�<�>jv�F�Ꝫ���3�w�����gp0љ��N��Nn�ĤܤKQ�	�VM�l�t��u���|���M��V<�j�S�7��̙O+��X�~��N�g��;��~u��N����}��6����r����N˖<�H�{ާ|�>ab��%oo>�M�t������x>��4�uq(,�J)�2ҋ��:�jN��C�;I���i�nÜFa�����q5�-Z�@�����M��/`1���{����zs|v���*�nq�R
d�e���
h��,^ю�y��oC�sӟ�ʲ���퐍>iq|5`������{����j�[<�3���{蹃b\�[t-��e��q]�:�٪r9��U+9��5�ye"��#"I��,�0�1,)��R�*�ό�s�t�&����7��Y힃����[^Hh�֑h��R�@x4od���[؇�<�^x5�:��_-3�B[d�}���-�=>	�Y|K��R������}{��"=�;���^+�_���L2������͡�NÆ7��=��+������h{8��C�r燙�=�k���j�Y�Q���Ӊi��:n�3�u������q��@G��ց���s���R�郰��ei�u��p�=�=w'���c����g�gљ62V�w)������}t�+�Z���4��<w򃟶�O�������V��E���ȸ2�{�^���o�\}۳vϯ]��,7��]�w��7"ۧ�=�燆"���|u�+79��垽���k-�;����"wa>�|��K�8n����$�wLh�vq��N��~B�'ޙ��
�M�h�@�cm��wP󣟐��V�d�&��]�����C�P�oO|�^Λ�E���2[���j�or�\�^K!��=
Nm��\��l�j:v�?i��v�3l���3V5�����{��d�#�z$��GX�zx��m	��{���w�=�ƕ�'��}�uz{�;}��Zf�5��NU����
��l�\?�$��lL����5�L�#nL/�J��-�n_lM�v�"�^�{�md�}��Ыj��s���.� k��;�z7��'��q�)�k>���\�⊁3���Ѷjг��#�=���c5$�s�1&浯�O�����PQT1�7'���~��ӟ����~�z�~[��p�����8zo+���D��B��;Km�T�4�M3)u�J4�)V����֚gRU�bk���Ml�����՛�RiQe�;f�:�8�)HG��UŅ�Kw�U�J�c���ד�n֔&n+�	muh��T�ˣU�M(�[um(i��ۆ�ŠXk�,r⛴��%�L�F��ZT[3p7v��6�V�kݩ�����b1��h�[�2�9Y�-���m�Dl�R��B�
�u[X�H�K�[��;l����Ҏ��� �KwQȺR�֯!6	����2�:�Tl`a�$��*�ST�FP�
��;V׮��ٗ�U3յc���ԋ.]�ԏ8q������P�M���z�k9,t�>!��>�ٽ�y�".�s{�/�FF�t��PБ��^`���z��<gm��V� ��q8ƀ��	X��+��8�v
�x��ҬƂo �]���E�ԥ׶ܪ�f56'�s4�Q��y�q�K�zi���� h��%�����*n�A�煥�p��m�yo�>��3߳=��m��6ucݭ�Ez*٪��3<M��E+o��y���٤�ú�M�� �-;zu^f��"�Y����/}��6A:��X���E&�lu&��)is�`a�n��	�2VU� ),\0�]��,���9��^����@��p�Y1fKU��6K�*˴LŘ7� M<k|x\OGS9� &�O��'��-�/@c�Y��������E�z��#m�3�a���(ǟ�}�ϓ3;�:r�ε̫s�˪F{�������}ߓ��A�s��Px��:7��=�����zM�Z�`�5��8��DY�MH@v�!�O�ӘPT������0`���E�B.��Š��h5�3������l%���Bͦ��t�p��e�&1�5�v,3-��ud@���3��޳A��D:�3;jӍqܻ�7�%�x��95�J���s"��3��"q�&�IG)M�U�AQhQid�e٭��sŷ즃�0 ��%m�Z2�M���	Ȓ��,c�!5u�k�
SI��]4�j��.���F>�9���v�0���Y���/sCN�]�
��m��˺����g9�&��GLȋM#%F��Dg��R�g��z)�z=�4�$�d�铧[5����w^Ҟ�K�d���~u�o��Ӏ����Eb�h��f\Ś)�6�1���ܘ�]O���_$���c�C���v#%�0Z��A�����vw�i��3���0��GE��l��cU��Fc@�P�ih��إ5���l˰Ǜ2WKr�E�Z�k@�uװ[+J>UPQDAZ���a�^
�9��&�O),���pa����<O���nb���p8!��݀�g�t�֊��tؠ j���H�s��NI=��8�~�K�Ĩ]H�ZQ�H�QJ)�ܝ����P�{��t�Ǫ����]>��t����:�H"����"��ﮱ/3�?osd�(ê��8�Y��E����._j�'f���磖�m�P6Ɓ.����ƻR�fZ.q?~#>q/���س�,��O�U��z2R�rv�P��
f�wXU'�St�N��R�:�5�T��" ���*�']M��:�0�V©1�nӚ�8,��~�R�mob��T�d�1�f�N�(�,"��l#Z�J�n��<
����Cױ��p]�P;�9�TL̹����^w!�*�헽��U���-.�УB�����鏰����
��]I�7��즨jPr"���h)���K������	?vd�f8�Lm�|y��VlF�s^� 8�,�f�g���3�fi��vzu��
���,8���JӳJZ�A>PA�]�v�sF�#q`���Lk5uc�u�f"B1��s�J��L�nĤ�0������L��a�f}�-�x��.�|��Ke��g[B�i�\U"�5�9��(��_?^:����ߩ۵���p�:� ��;Ɨu^ʷ�����S�</El�d�+����PV�fj��$qrG�j�h�'���{���3���{���9ωQ����6��������s���j��("4�\޳q��]K��� �B�A'� !�a�v�u�t7VxPS�d@��cL��M�X�n�s)0b��TB��In�KIw;*���<��V�.��^���c=;�<d��X�j�b��7A�����Q���b� �͘ū��O�~ݴhP�q���t�n.��7V���n��p�����RE)g4a��;��z�=�M۹Y��۾��s��u;�y�������l��}��xNT�֜�~F��_~d�78r˵~��.;����6�_������U�O����|�C&|5P��J[�g����r�i�ȯ��q�)��8g3�Z��
x�,b,�p'|�Ś_r��%�c6�e>k�f��9X����15A���|`�|�;Þ
�j�úuy싼�s;�I�I�8�cw �_�7���\��)��{ݍ?Z���]�`�����"c^){ �`#���#	�:������5O�^�
���o$����-�W��c���n�3N{��{�6^cU8:{����g�'��6<��RrJP��b�n)���G�qsϐ�|72v�d�І;��:����_c^����|���LD�PG&>�g=�������"�*"�"5�o%^�[T��g��e�H��A���D�U�l��Rk�װ�ѧ�}CX��U���ww�<�}o���c	]�Z�-��x��MQ��ܕmP�C�Yҷ
�W"�ܜ���5C�i���҂Һ��fU��L����9Sޖ���a�@tǞϹw/־���J5�V�
x�l�I��s0���*r"������sm�(�*)H�(����Ud<��#��@�����G�����:Xmb"�0�;1�}N�,�����!U�wsĹ�����M��� z�nh��4WZ*������U{~�J>(C��Eu�0SU���>��1���XP��7��Dj���#��hs�z"_��0�]���E�}{}�9��u���"���11��J��b�Lc[pMqE1���*
9�����6�e���0�0m���Wd�,.��Y���Q ��'䷭�m�}ݥ��xxOEt[q�9�ʷ!���)�@�U�F��C�a(~aB��M���`h�\��j��V�-P�ҲIV������FZ�U�C�U}B9�Qi_4F��K=��3���h�P�ک��W[�:뾼;y���wp��ζy���_�CF:��.�i��b�4��4J�T@�%ZP�� G�( ��s<#�����*�Cn;���e�ekǙ��.iݔ���q�í����i�QV��EE=Ee
Z�A��!o=�O�.����Sy�}@�+�+���1���^#���u��[h�pJ�����sZ��x�����1�g
�4+U^���F.��%YW��YGJ��O/I���2�S��J��D����|�n+-P��J#Yh"WP9��uA�k���9�c0"� ����wnf�.\��{W��6��1}�/\@JiiV�_UW}w\j���~7�e�^ 4[A�ʶ�|U%G�@-�?_��i��mJ�5B�h#U�SY#$�|������-R)�z��@0нD x�0�{���y��5���\f@S�Ұ�;�V�̪�DϺl��h4��J-(֥[G
@=r�S�j����Q�7B �^s�%�H�1��FR`gy��[���9��l4g~�c:�ڨЪ*�H�4�����.v����Ϻ��kMQ��B��
0��(R��7X{�����}�ؚ��*�6�Q�˛�f��3���eUe
�!ʤ���T)�o~Ç4J��n�vQ�@�>�+UHQ��~���3Fr�Fd�����{҂Ҳ��{o��.�J��j�d��R�Һ�4�sR�����|���kޅ�A �E�{2��7x%��hnb���]֍ȸi� �{�9�n��{����;�p�v�I�.a�.����h�dv��b��
]����-֫��l�B1��2[��2��\�9%ݎ�k P����{�6��Ye�,�d��<�2ت��4Ux��/��~!V�kR��'.��SE�vZR}��g\єn�(�[����%J�H��7/s5���F����9���t�p��"�|<�jY�s5{��m�w�$߁��;�(_9[��}(x=g]SK���t���{��!�㱚R#�� }�9%�t�)�Gni.u<�r*n~#�9��A���r�����DV���fn��Y�[@p �r#����=��}!�@�g��q�o=R�^��f1���͞�I9at���ǟ�/���k��ajY������
��q���v�axx1�f�m\�`�< s6�Ԙ�B�����
�.bO%ͯ˦گ���aSXy�j����Z�!Q:��\�H��@j1ZDUW�zc�]�Χsxdg���v��s�/_��'f�<Q�v�;߬ߛ~��|=���(��Sb�a뻧��c�y~�o�~����	���v;&w�<F��̳(�5x<�s��qlҕ��yl�K��Lb/�����3��틎�-I���\��7��{���AJEiUTQ�PwY�{\�.�y_�������|��{(^����h�ji���8���	�4�j�0�NyH�h�l�r�\{��@�ߵ���쎳U{'5w���Fɟ�B����}���4xc#"tP��'�� }�2��c怮m�G��3��-��AA�R��[2��F���	x�I� ]\C9n�dӞ]xX�TI���ݾÿ{Q���(U��ǯ��v�\pd3QZA�~��)�=�F�=G*��;��Ǜ��.�3��Db�ww�n����4���e#Ϗ��JNI�X�hx;�-S�T�!Ο~��+��P�y�/Z�K[��7Nwu��^5��?��o�Ǽ���i����2��E���͂0��`��=�Ood�	�:20
���gˢ�Gx=� ��v�j�b=x��^�
Zq��|HŹc��,s��rq�Xv����7��Q�k=�6.W&�"�M�HI��\�X
E�+�
f���(+b�Qˋ11q��QbLƲ�`ba-�&��dk���B�׵��Lэz����䶴�������p��	�Һ��6�\H�P�S3eZ;*��eͣeMe1R�#t�ۿ��x�V��1�wZc���# d�#6���Թ˖���\p̙�t�ˣ�B�%���jM��r6SXjf�R�m�q5�R��5�fa�����LЮki�\�94I^�3Q!�u��v��J�-�X��;Wg�X�*���דK��C1#v0�Q0�fؖ�nqshF����-�w3����5vX��u�q���j�Rh�f���lΎ���Y��ԗ%ՎJ=B�XM�8 Ȥo��$��-��R����| �!�4>6R9x�7���֢��5�b�0�`�����a��1�/C'��9�My��MƵ������|n-̙s^�i����m����W �OsN�1�{���zi̺��d���8O�>O'���j��,���6L����+��ۧҜ�]��p	6,6燽ӹ��7����k�a��<q�g���i���e��z3͵�n���c�� z��Y��q�{=�s�*�^<�:[
:�LPiMSQR)�������cZ��^ui�����n���u$è(F�д�6� Z��4��e�ت��H� �%�9qf0^˘�BX�����'G�F�'�66���{��Rs�Y��ֽ'���]��� 6_W;��f")��p<:��#{#��y���Nd�&
&�v�}����}w����/�-���z��a��4Y�ıy�!�v��f7�;}� ;L�G*�vwu��u��㺛I�ݚ%��l��`�9l1ӭ5 f��yx�	$y�P��NI��Q1��rb^/Z}�j�Q�b���Lgѝ�����\ԏqw�/zm۸�Lb:�� ��Ӓ� ���Sש��:�h��WMԓ���)�3��¦�<�y�K1�<5b`�$�xa.H۴ @�s��s�c4�3���v���-�l%�3��6i�Z��f���5�q�]Z����iQT=@_ܻQ����=��q�n�z�;�E4:j	`�k1����Ԏ_ÄMvf:&&XgT������s�܍k4%���y��l��`A�/ sY�U ;�Jၦ{�Sa�H$�S���$<k1��%�ݣqFS������)�&�v�
�oL	$�QTR�O:Ž���b֔{T�T_1��ܓ��~d1��,pb	Ap�;��ϔ����{(_>?'^�ʍ��I�kO��R��x�䘚�*��������sY��<<���i��靧_PJ
����]憨��]��v3�2�W���((�J���cy;�y�3��ϻN۳��2�dCRָm��.��Qt�;QsV��d�+h\0-��n�f����)|�����u�{R�.�m[7l�S1���`�ڭ�su�:�z��,�:�m�����˶�.(��]�,����ne�=���s�k�%PG���?�Ͷ�L��j�é3%�� O�\ɞT��5<��R�{�B�����똑�n�D�����1�=c��7�?iY�7���TH��(���ٵ̽UVL�2�s<�,{�eV�tk��.d���N
��,ˌ=�!
W>��	�6.�*Т��4()��&d:��(0�˾�3�]�g�AD��ɍ�,��5�!A�#�ݨ�h+Y������px�=l�&�c c��`"eZL&ؑ��O$��<�����>��1ǿza�����7��U�,�O�]v�B[�p��g�*�4�����;1��q��3% *�T->*�1��o׉n/���;�i�&hj�>{�>�8Ó��%a������}8��[�:+5m]V�����k�|�M+ag�$�����=e�x�^��q 0z�[/�E���y�:��+�3����1	�<�ۄ�}�;%�D�c��z��^�I�{���>�4�MRҔ��dTU5c;'s��IU�N�>�����e�Jv��7��g���j�C0�����K�Շ����|�(J+F�o��Q�Tu���y}���IA�L�w3T5U�^��/ZWu�5�"W�p'����K�.����YBn`.�����)�d@.���GTp�z���Xl`LXٳ�
�]Y�u�٢�a��V6��j幡�b�1i��)��4�r"����BV�D�Һ��r��:y����1��<�m#�l|�&����5�c�ފ�Þ=Ǧ��bt�S��PV���DH�ˊ9,�R�@>�[=�0��n�4��r9�N���-c��t�qi�I���v��~�|x+�bEI��#m�$�y��KLO7���x���Mk��׸�T�-�R�K^��j8�ۮQ(�y��7��vQ��3v��zb��3�4��$�1�G�/�3��~>al*��}峣����,kU��`!������co;|��:�h�ƴ���I�c�:�{�F�K���#�E]v�I[��y��Z�ي��2*��;cRO=2�U�[�e�{�u/�9�^�t_�u����$Ll:�r�Z�*�TkJfQ1e�&V����Mȝ��Qa��쎋��v?k�
��m=wt�u ro�v���p|���O��w�L��������e8��"<�>���.)�P�yB�y�;w�8g�{W����������x���s�~�cݼ��|WEҝ�,ݬ�g{��Yˣ)��`덕e$��;������exz���w�i��[�oqM�g",>v�6���r�M���#x<����*��Z%��+��|L���>Oӛg�]&���[���\�N�~�g����֗AT��(k;����B��~�-gY�#��L�������U��!�^�˽�
�Ս�ѧ��Iz�2����`�8�(j���3�uj���47���c�t�;A�Ji�ipo�CN��;0���7 ֯�
��f�!`�q�Ϗ{�;�X���;7c�9;ޘ�����n�n�`�c��3|��6�����*4����$%��zv:Q�3&�y��/e	k�@���c1�&�@��l r���J=L�1��']����\�� �m������O�	�f5L�� n�V9���l��iJݚ@xyo
�2H.���G��K1}:��&�> =������Sf.;���N^0uȺ�b��i�y����;��y����z���Њ�*ר��s�q�g�½
�O��2q�3�%��s��T�4��tT��x�wfvx�B�0�kd�XN�Ow�aF_c����P��L�����l�`��f5��zͻ����r$	�x�]�#i`���\Q�B�k���o��T�:�P�
��𚻗�ɑy̼w���0=��6[��W\�)c�M���m,��#��3([e�(�5�X�^�-9�t���M�L����b2X��j��Ҕ��"��ͼɃ��2�"�Dpw������B�x`W+�Rn~�� �q���@�P/�bxC���~��,Rk�ފ�}#���*N��r�h��t�(fՏv�ۻ'PrR,�w.]�	��x� ��p^OrN�( |�}`�|�u%{t�����	w��33���S����EY ��"��I���PD��zG���U���U��?�����zD������c�G��f1G_����͞����[��z'���>�sT�e�p�`D=N�c'MPx�P���0����h�|gvp��6�<���� �-�=�;��ܮW=&�+�@��T�^)]��Ȓ٧9��Ǽ�Y%�!(ZUU�E;�z1��x�\��L��x^.��m����>hG,� m�\�=�V�Z��4M�r>o�ȝ�-�������f��Wg�xx#R��p�<@��Ҕ{�;��<�f2����/����r�C�K�5��64��{��9L��U�	��4m�I
&�*�_0Q�R��U\��=֖)4v���{�K�6)�k.9�ٜj�cJ�u�NK�3��Ͼ:��9E�Pq1��z_��p�(���9��~�����w��&����?+��-H��/�xyn3�n�j ���c����d�`#�D�(�3O��v5�ev����lV<(܊}9XЈf��2xz���L\��u�A�J�k�-iV�menl�k�p�a�-b�X��j�� ����sf6���|��[m���e�Y,�[l|��F��6��fX�� ^\g3^{��f���	@� ��*Mx����[,��3l�8����t���EР���
;/��k�QA�b���f�ePT�X��X>k5�����;,��;�Drlb�,6�S71�Q��;�"�����m"�a��9��Պ�sm���!����y&e�Nh��ҭ�s0G����X��$EU �4��'��w˿j�Y��MQS�=ǘ֞ ������qF�҄{�, | �p�,ǒ���`�_P��'�8�)�s6�7���tB��H��n�у�E�$]���'
5&trO2{��`a�wg�f��s������"���1ntE"&�*1������EF�JZQw]��<���{��o��k]j���p�)���[�{=xr�볞�v�f�f4=6h���������A�B&�Bmy�����}�2C�f1GS�2Mm�yǪ]�%�y�m��<r�W�}�ܶU�Kc:ww����c��oL��E�(=R�z�U�.{���m�4¨�����,�%R�IR� ��D�86u��qN�d�n� e;t���������ԣFW&⻂ıa9�Ɗ�Y��z:ͧuK�ՙ>a���lX�n/U�B��.e9��#��Oi�H#�(EG�jZǁ s#�Ah<�雚�K�y�nU/4���_�v�
�~ۏ`�Y�.��`�G�����x�v6�Ox�w�X#cn�޿�KR8.�D@��3PS�SM9�P`��:�*��y3hM׆�I�c�D-���j����o�{5�n��ͽ)<�����L��8��CU3Sn���K���wX�ш3p�a{��v)޽�g�W���px�6GXT�l\�a5Ï"Ӱ9Y\�B�He�M"q�{�n��/C
9��.�ȹٜ��=�p����pm�>��tu��T.�0cxt���](,��R��j���4�r�-�,�b���	,�i^��3�]��3N(@�e����t��:�J�Z�*�ⅻCKu�:��c5�6����[̵M���\J�k�[Qlؔ�6�E�M)G�� g"���M�ҕ�KK-���1*��U(dF9#��Tfn#G"i@��Q�B	t\tvss2����٨٬�\hæ&)J�qe��J�G9m��f��"�.-�m��l��0�P��b�6e����.�rW6͝a��)\Sq]%��L���^] .�6���P��4�r���J���B�R2��&��e#����+�i����_P���������.��K+@~\]�ݱ��*�v s^͙��e0x�֔$KŁ�% ��[�i��ݜ�g�����o���4̠��e.C���!X['AR� ��L]��,��%�6<��o�m�o���_kG����듄�0�Y"�ulj>=���<|q7}�X�x��&���z����a{��wܲw�+r�%��������<ǎ3nN�����gzݝ�|�/����%��)�����M�ʈ뜮qt�.��]�8��.��五��#XY�MD�Х��ɂ�F�:��K�8`���U��ZX�#"QQ��9ue���1l�1c���p����'�8
1�{��rY�y�My}0Pq�Aj�PP��'};�$+�:9'�0���,�G�8�v󱒁�f�2�#���g�9੸��>￮����l�T��l���K9z���� zx�3̞F�[/�^����_9q��ȣt�1�A�	�"���J�I*8��ԿMf|8�����q��W$i�}����6 \X̰`I��}�t����
`���q1�y����]tS4 [�h͛�U�~eٵX�"C�=��7� ����`y)��i;��H���ɥ�X�ksh�,�J��O��N������#"�**������]���Ͷ��A��ڝvh�c�.�<���-�j�B|#lG�]�V�B�i�gLj�^����<����W��'@+ 
)ؓn�<��3A�!C��26Q�1�y��H��e��y����,iK��N���Z"!��ZC��wgp�u͍cN�D�H�E��B"�I�F��?�?Iғ�_-�:�}�~�|khk����9(�*b��Y�m#)X%>%��g0k� 9��Y�( ��5l�'�N����혽~NZ/��w��%>B�'۾gwy����R�L`,��-7&!�ܴpº^Bȍ4��T̈́`���־��/�"�M��Ь-hŲ�i`Dڌt��̱��כ��4�a����\�x�JjS[a+vֹ���9͔��씵$��Ƣ���J�	01�Q�vY��dÛH�P�Ԍ��|�e�]��2w f�f�fG���{��u��5���K2y J�7TS�LU"��9�И��䦃7:��R�V̹�>|ߗ|��߽<�TGXi�$�|��Y�Ǜ���ܗ�~���������!*$djYH��D������~�{�9���_��Y���={��\`�3�x��~z��'O߶����.��j�:̨Vr˦�}L{�������%<�Wu4�{�y1;sL�,��1�`j���>T�12��U���R5#6��Rв�"�ȌU���}1x�1�Ҫ�g@X�:G��T�b��'I��k�'�m��|�����w7+U3��UU����������������A7����&TZ�����Ԟ�i�l�w$�\�D�f0Q��I�]/��nD��*%�pd�qY��V&���ǟ��q1����VŔF
B�����0T�Y{~sz�ͽ��ֹ˷�@��a����@�R =���B��EӬ0h�F��w<��{��)�k<Z�<Q�̹Rs��4�5��.��[�f��ƒ=�� [��M0dY��@:�(���'^k��\iQ{T�w4���zu��mv��0��A�b�d�iK��[��!,�W����\��oMaU�#L[�w\�*f���1���Q�l3��rV*��}D�2����u�X��LL������S�I���5Kd.0���q�G�r4�G�+U�����	����8�s൑�f�f�f=<Uc̞Ag�vc��iz����	���4�k����&�I�&����;;���\Tut�]1u��6�ъVσq6��(˵^ �Z�1I�		$EVAFo�j��o�g��a���>��7�;����s���G�7<�0׃C^!x��翷�{� ��+��Ƴ5��V�$��x���t�T��7��WL�L���eRz��*KDlB�����f�d �.j8�A$d;VK�d���e����G�8L�p<Y,�� ��Y�=��F{#��4n������<��;Rz�_�10��DTQS(�äBi~�0���l����s9��ۑl����J��	�VE����;n���lCnv0SUl�!�ٗh�y�`7.�b��y���� ��_i�'c�z�<�}�tI���]܄{���f#I�6���j^P%�<�G���^��3�3�sf��_�Z;i����O!�bӪ�*���!�O�@�׹��i�PH~��Y���sg
���a�9����t���z�1Yۥ]��탩�*�g1�������2�˼3�P��j6���_�N��3zt�ܢw{�������3܃Ģ�垞����p��x7Ϙg�%�+^���|*�,�u��'0=W���ox;�x��I��,(/�7�n���h�}�Mڭ1&����B�)x����������nnLs<��..rjb�E�#J(1�D������cH��Qkx�7�'���p��o=_�}�s����K�x�K���3U�8!\塑(����!��|�����	<����y��I��Ykc��G$\����Y��Jxx�� �C*�z�F1���b�9kT�WG/p�s+_��"�$jBQ$1�!$TDUB����}4�ފl�����-C�g�J�4���(�������Ǉ�����05J�h��>N�3�kEx>�)�Xvr(�H���/Lm��c5g�P�B���ya�tO��~���F/%���b����+����i�D������7ҩ@�%�c#qM�ɑ�Z3ZZUlM�ub�ҒŐe�)-5��ղ�.R�U�c�Жl�o�ݦ�ےRIJ,iY ��U�d �!�9���k�R]�xc��n��ƞX��~��������ڧ<�~R��
����Ps9�Ե����I�2�����V����y�W<u�g������Qڵ��2M.�<���!�ww��q��v(��0���{W�s���N��3Y����e��ʈ�SJ(F0e1�A�)a�>%B(�IrGJ�x��7�I�Os5K6 �čs[�+Ù�s���Y�ݖ�%�d���OiG�~Z��9.��0��1�q��G^��-���dw$�Ӊ�I�M	(ݴ��N�'I����eĴ��A�f�l��i���'ڼ!H��RIi���e-))�RF��/�1w�g��ם�o*�K?M� ���g�j-�(ǃ�§��kZk]��]�������4�f9ఱ"x��c��e#��o+�߰�bI��%�G�����1A�W��v7LК���GN9��6"��V��|�\�u�d��i�a�2b��A�����a)������۩1�O��{m�Ù'���E{-f�ږ�*S;31v�N�}�����)�i���EҀ�e�G�x�S�-dh��#G�,xV��G��Fy���cR����f9���
[���Q�k`=s" �+m��������^Xy��1��Mh�&�@V�`T�Л\��ա-4#v^�1d���l0����5�pR�t84ZZD�rM��Y�L���7�qB�)l),d"����V3��/7& ��ţ�����6����-��г�H��`�6:�w~�hJ�I=X��$�N��4�����4P�s�$H�����t��'�8��3!�{�aH(k�[Q��]��jb��eQ,WX��'�{2�;�V��O3�<�M�_n�����N�5�5 �$����J�г���3v�}E��W�v1��`�
�n�;�'u3��rl�\��c�uX��4��R��͐�v���/��iV�	��uC h�U�¢���$y���y�y�]��x7�C�A⋮zZ�4nl8O>���i���K<#6���{0��|u�IY*�B$bH� �{�������LщqD�[���Ƅo�+�=���U�������8b�ˢ��; �VV��}|�B�uw��ov���+�Y�zٷ�J�&
�i��n�s�E�?s�If=$�i�3��YS,Ǌ�5wO��#�[H�uʾ���5��oY�q����u`BTbI�"� EF����DEI�E0#���;�ܝ(�*<⨮nE˱0�Jŀ�x��k��~�]�߻�;�4r8���
��
�f8T�Tl�:e2{��ٰ{�ܝ(��-s�󹒋�ʭ۬��I�L��VCB�E���������u:�����YH�1�	��s*����M�Q�r�i��G��!�!�������v�Я�;ߗ���vU
�"ݞ:�K��G��YbǺz�)��z@�&-m�����!���-����(����m�(3��m6��ނ%����J�6T`�)n��/����Ǧw��zN]u�y���z-��չ!Q���GZ���G5�۞�M ��7��i�y��w6׺N�j�IR,k���au���H�_�1�qT�����p��{��7��`ݷ���=�O<�fУ��NM�8-�,�l���S&+#hgp��Zh�t�0R�B�]����h����PuCqL+n��n�a`�0�33h^�t�YK�k� ��1�J[������4��0:���m��5ĲYzˆ�n�2�+)s�n�Y�\� b�B1Ee���55[T�d�@�	Y���6و��+�bKq���vöыv�0pբBa@�f�����y���!����`�s�e�ƶ�q(��(�4�b����(�k�^,�X]H�cu,h�����%�V��R*�f�E-��*�r$��CC.e��Ʈ����WJr�;��a���6�q�d�m�\�`Ҳm�5�����=�x�����y��ur4)C#4�!;����P��ۑv,ۏ�����t�=��QоlL�Qnx���>1���^�<2S0?�9��'�]�Q)=c�x����C4���n�ۥ?g��ڇ��0o/��:���1�|׏�}�S�gy���k�{���w�;}�ݸ;{գ�J�m�<����#IH^5��d�3�h����l�d�&(��Zi�*1A���Hh�L�h�j3+Z����˥�K�v�äXG%���SV�Gbؠ�����s3AJYX$��7��/�-*(��F +R-(F%]5���n����`�H���.Y�3�.��"a]��l��2�(��� M�!�ˉ�]�o(t+��!�q9#�����${��n3��r�4�<�}���:��7��1��q\a��cFlͣ�w��_�q���Α,x;�7�A�oF�E麆؞�����k:��w��LrB-4��H�I$UUU)%-"*�1iJ�
K���I����%�g���8(A��؎�pg1�+dDS7s5�r:���0d�=�s�Hǆ�L�˺+Ul��4�W �����z�-�py����o'g/2x� (d{���8>1�w�<Q.Cݸ����. �Y�.#呒vn��m��|I@/"H�L�PZA��H��ZDQ)h���Y��c�b\�@�믧p��j�@����=*J BN&�� �v�&ƛ0&����޲dd���3e���铘4���K7s0�f��7Pd�QL�3H�=r���7��Y���5�,�r4�z��b�c�R>�m�W�%*5QH��H�d�H$d�H�Q��) J)
!rb����3���c���V�::����uJٌgKt�
,��$�$�D�[��B#6'G�'�C�[7K1M �奏x�O
��B�u�JGx���H�P=x������-ܭ�̽_KeN��E�Ʊ�&�ఙ�9�.b��������!�2Ev�E��8]��FmVh��;5 �K[�8e�Fd�,]v���Aش�JE�JDM�n��%�ژ����Ki@h��0d`�"H$�D�F)!am/]tץ��b��$��D���N砉��w���x�.�og�a>��淓�������[��d�gx�x������3���zm��Χ�q��r˅tr��p`�����'���Z�3�����Og��˻�=�&k�b")���ܿL��6^������;�LdBH��iE#��,R,�"Oa1s~�W�m�<Y5���d.�9N���u�����B��ww�垹a�c��<i6:g%%bZ�0m����l��������[�I�q�0���
����%N��/� ���*��M��"�
���Z����m����"��! �`������J$�AIH�-�� ��A�u�8։N`���P��R�#�^)���I�.�$��	b�kR5��0}{�������7I��b�| <�����/�Y'�P���M�k����b���*�����������٭��5ܗ@$�B��� � ��(��JH�H�2F�JR	/�$����EYvw��o����OO�>��X��0��B�Ѫ���/+^�Y".gh��4R����cy'g1�����f.��,�,zЪ]�|2wa�e}ְ	��NEG�j=˶���,,�N��s��SNFaf�E��1�Fܤ
V��8)lt[[�#�=����2\ej��Gq��s��f=b��k]��C�1&Tb2T�,j+j	H1�VE�i�9�c&.��w���q�8wp��3��:��tz�4����\�z�rG���U�RhD=y��b��8*���r�\�@��c���%���='��۷��bfj�líB�T�&�z���DpV���O4T��t�4]Tt&���ʆS���@�F�"D��RB@�EB)%B��Ų��{���3n(�~�sA
N�d����L!�|v�o'w]��ܷ�}����`�r�-U*W-WQ��#�؆k	�d�����y����<�xDͱ0�)�u(3�Z-�6l��^�&�7iɇcd�lzǊ��`�r��E��yu�@7�F.�z��PG�zj���U�D�Q\���Y��:����kc�g�}�X���l�HiA�`���3mT_�3�;Mº������V*nF��}TG�\��1?B�gso��>�ZOy��\[lҴ|��Z��q�O[w���~���ߟ�{�e�I�fݩ��H>��/�O���{�3���OP+����|?d�5��#����C�ʃ��������c���(*Q���y_Av�mS)�"#���,��}�{x�b���k��1��yO%�vvv�xv%������t����8���қf�|���{Q%.[�T_�hcc�C�r�����:$�Y0w<1b(��?}��U�g 5�0<���M�t���Q�1��)���⡤�w��X�)r�Ӓ��w����0+�yQ�:���8�iÞ{�|���w�����]��}������H�"�J��Qb�"��%FU�|����x]u����\u<�0c[�Z��(9����+�1����û��Lb#������>І�g�'�[=kW�ݨZ�Ӕ�G��Vn�V1���Qzs+]5Q�Ś���ψ9�j,��! ň�I �;#``[���V�?���'	�r��e���D�"m��{���}���)'���Us�4Q�UCE{��ӡ�av�=�eq�<8��t�u����\�˭���[�"��֘v;�N��{����g�.�4�\ṫ��4����,��y�h�a�u�,�v�n�ZTl���jk,0��T-3�r����$&��@-8 ����t�z�;�:�J�UF9X��/|��C�8�wx�`���@#��wM 5��6�L�7���k����a��9��O%^"�{�i�ƍu��ګ��{�v�譤�@�j����Лס��2���g�[}x��EI%Ac H����PT����x�@��a�ʇ!P�I���rr;�J_R�r�G�އk�fd����z�fhkn�`L�e�qe�'�ܤ�g�z��3�冒�]Ǽ۶����m�p�v;{/(]�Se+��k#�#�HI	"HB	$�B'��U4�ή�8g���-��.�W���2|=y��b�s�Zj1] �-e��O�=���8��Їr��3a����^l��<v�{��e��]
���� ���KT�"��ʻuNcdg�\�19��qRE 2A����%DP�!��5NѺ�{��H�T �������Yb�1����Ğ}���s�]���,�(��i�P ;����֞Ux�9΋�]�(r�CL{�T-�z�3�r�CMkO�o��D��9�h,N�[Y���jq�� فj��	���P
��+�
2�2�D����AR`+��k���q�[)m����k�`A�ʗa��mL�f�Œ�.�������ke⯐�H� ��.�Pv��>��{��};�������Bd z�Hng���xB{�%�E���P=V�:
���(�������w?>��}��R�v�c��dX<��bxO�A�2O��)�Y�\�a���ƙfV�Њa��e��5�GU��JZ��$��a�����<�9ܝ�<_'6 =��Y�2��@"!f�8�&��4�\�a��ޞ3�{�,W@L�[���2�<����5#��p�<�#�_�d��w>n��,��2�I��LEzn%�@�}�l{ػ��u�����a��;�Tu*5��	�@䇹�=,�gK��㖢���ÆX.�l.�N ݴx��3;2c(��(��R՞���<��ߒOo��n�ON(��ؠH��dxx��.><��+5�q��^��2ג����n��պ�_���y�k�F�AiE�!%�$�x�;$���]�����������&#��A�����N3��It`��I��=� O	�%W�����v;W�-Mks'p�@W0�C�W����r�;�q�x[ɭKcċї.Wc�(	��.�C���9�+/g�`�yl[�}[a*@�Qw�}��↪W�7yM��^�������s���)L'SB�lME�lU���6���ǻ��#�T=4���tf�����-����8�$���g���Iz��V��ևP���VaȆ8b���BҒ�PaxU��u�jxxt=mV{��t�+�LE`�:�W�d��T�����Хr̫=췋�L�K��v�~����o�.!�%�k-�f�d�b)���.�v"����[�Ѵa �sc{Xb�r��1�*X;kpR
]f�K��]KJ�H(�͍�5����Ҏ�ݒ��D45��Gv�#u���fh1����ue����W6�cm\/F:�tqf��c������"�(̥��\���ɥ�s�-�Ֆ:닢�4k���P�,`�0��ź�`]i�k�m��ZQ��m"�lK1���,�Ml)L���U1t���!a�[�e���#`�]�g1D0���;mB��FcXk�J?���|�+rRn)��%9�M�,ZT^:�hk���Ь���]t��8�� �<<TXF���l�Sk�T�A��j�u�i���������n��龐Xh�Kc�R�N��d&���M!�6{��뉡(� [�$���s��+#�t+�r>O�U�Ǘ�����E�Eҷ2~�>��OK(��>���/e4ֆ䚉�_^�n �y�7�����Ú��������g�ҵ��s�oA^!r�Y*d��u,e<���8b.�Y9^�G���JU��8yoO��9�z/���3�݄�	��#D�v���9!=�}=ݞ��n�;\ݶ�Q���&�l�.�`0�,�γ]�kV����We��m�[	LUh���-�4k��G	`co�ũ#R ČDP�DddP�E�J֜0f�%�0ܤ[�.�	�S/�>o<߯��.g�|<og��l�YA�D��sjH���}E����q���R �a�2ͼ{�`��G+"FŎff�Rw�p�d�&E��0A�w��.���o�1�+�mS�H{v�d�\Sk� ԡj��BP�b��#"�xߦ={�'��$��#�������~h�5��u�z�*ԁXw���9,��I��e]�tæ���u��7���G�N��ӱ���)t+u ��]��ۉ�E3�i:���״����[ˆ��q��ڵ��}�9Y!$EM*�a$bI#�ZT8X'�즘ZD��5���<W,���w�y'�S��}���W-�W:�9gt����� �D�v���Y<�o���<+���\2O;9���ڏ��,�J�������LXS3A�e�CS�����Q��r̠���H�R҂�|�{��n��~OQ��M�sA|�7�b�MYD�.H��l�w�n(���5�ÆH���~�D!���<�x������ӎ�Ms<X �nǽs�Lp-]��y�;:g�=i��;&/]C(V;P�ֱ�DH����P�-�F3v`b�a��(bцٚ2�$�,��sn*�B�ؐ鱅-�&%�b���Ulں��h=����]�e�,���T�M�6�vp�\2,����Z�Vs�� ��`��԰k��#��C��a4 g4�z�0/�qD.��O\��������Ǹu��(GKRԩt�2���~���MK�w���U	1<༿sO��U���ث[o�e��z����T
��@�I���@�,����(D���y9�vC03��>�2��o�<�9���%��:���}_�|�[��Y�\Fks�͝Uׯ|'}��y�߼�C�}����WJ�S�2ŧx��klzS��O�˨���uN�wv�e+Oy�j�,@���3��#H�����"��%c��;�f7T�nT=	�ܵ���^�~��~o]�|��}�tYn:ťB��.��a�h�ܜ�g�"S��1�~���4^�C�GZ��9�ڞ�T�g��[	���HT[Bv�g�}L�;o�ٙ�[�9 ��H3^9�I�9��� �ѫ	��P�fA˻������L�,�t9vSeP�ü�O`�=Q��<'�3eӴ �@l���srw���B
/�`��m��_��l�/�UDUg3Nx�떪9B(u3���o~�|F7��n�j:��koV:�e�Zl�"�Z�XmJ��.��Y�b\��ZT��۶ٛYV6�v������%�UJ�����������WPfc����h�b�:�|�h��,�2�x.Qon�S��~}����Ja^����1�v��=?}K��z��jYV��*�Q��2�E�_K$��u�$K����x�[�2&Y��c��D;��'$@)�)+���p��u����O$�H��k�]Ή
x3���1^ns�X�΋��3�r	p��ħ/�!(���<1��O3@,�C�7��P��T��N��p�r�Y�"�Ԣx��c��"7�2��4����Dl�nj�'��
�������O$\�##��o�p7��o�dI/y%B��ط�nn��{��FN�-W+��bYڜx���b8t�y�.�f���9~ �1О�h$F慵�-D��i�+�������e��L��bG�_���%���P��m���7)͛Y= 3x��GC��\(��򓜡��׾��[ƥ�E�ܨ�����zd
{�K|�f�����o ��8R��0L��}�G.���w�����4�½�P���3ݤ�ҾZ��p��ͩ��Tu�KX��L��|�س�3:�����h�O<����f�����1Oo{q������}���9%�
={s�K�����u��U���FU�;X����o���ͫA��I�Ȕ�1M'��gmIR�!���y��vl����s�W��X��5:-�֟6{�����h'�0�ȶp�#�4S�> ��F@V����H��/���1�|�xE3�.nN�4��] �p$���;`⑍sE6*�C=��!`8oDI�aJ���u7h�U�Y�<e�6�ӭ������S����ܬeI�������A�k4]���h�V�o#�/Lh�ұ����5�r�j�哤Ӊ׶�|>�:���.6�tt,����A�6'�<�ǯ�.�u=�Ƹ�����]��`��$g4J�'���M�K<}ή��h�i��[�cg�*���v�}��D�����c��"�l�{��v]hR7kY[��7�v�l���B�R�IR�6 ��+ɱYK��wY�E�\Vj����t��%��l�8�y��l2����Rw`Ht�?I)���xtJ[�=מ� ��+T:�S��;����L!ܨxF���r˻�`;��{S����ǹuuFh��2���ܞZ7���3<vն6fN���7w7�Y���E��4�4������U�(��H��C�����[}0��ϫ���6�Lof6�]��$x�"=ܯ¥��:=݀�n�7�p����ܧ��	çy�@_�f�����<�w+����`�hf����҅l�ǵ�b��ʼ3�gfB��$�	�
-�	�Ɯ�t�Ǽ}�;�k�46����������p#X79U���`Pp�4@���J��g�4��L`xxK�ǻ��ysI.������Yϟq;@��U$��1�yu����0��h���@D��@%ɵ�&�k<W���$�������h����n�;.�g.� C.�����73@��)Ϝ3_y�39�,�����y��P� 7S�R�3�Y��0zV�b�x���e��hf�N�"��N2zîr�� Q�$3llI������#(��P�*��7&�Y����VV6ƽ�\7���۸�$ݵ�[΋��jRb5�-�2��*4��
@��W%ތB`�0Z�b���ߟ�ט��84�>̡i�k �	��m|1�/SB�x��L'�ŀ|Ά�C�R�Z�6 �g2=�|�<�Y��\Ғ̩4%2�`��wS��<s@�Ú$��:��Hk]�צ��w�ܹ�ؑ.����V���D���"2$��^'1м�ȕ�Hh�B$��l+�:.���xN`50��\�m,tR޳����N�hʴ�e@�&���O�?{��g���z�-+���4�73<�НlƢ�g
��am��޸�
#%��3FY�m�ܑ��R�Q@��Q1|�2gx�NU� ծ�Ty�<I�x�5a{���ҝ�4��f�.��h.�&��ٞg#�̅O����Jx��]i;�j�V ��8T�z�:�����Cs\;+����gj6vt��曪k��u1���`{3{�q��(�b���1��n��g���X��E����Ӥ.���
�R��.�~���~���T�g����.=��i-ќ����W=��Z�'`�5�`��/x�������Y�ͼ�m��e�P�8?=U�O�\������ܷg>WIӧ.\:t��nw^\���GY����+eK2\�q�lҶR�&�l�eT�Kd�i��V�b�R�EmI����M�V�F�[Dm"���U�Y�?^�����S��W`m-����j���&j��ʛBا^��m�'<��+am&ʶ��m�ͶCe�����ll���M�[lٰ�ڶ6��e�[#�m��ʥ�ʣ�8j��T�e$���
U��Mp�]*m�UK�G,KjSif���\dM.4��aU�`����,�[@碸�l�6+�&�mP�,¶+jVÆU84�YV�M�lV�[B�]��%��N�p9X���Ӂݯ���owB���HY�L><���}w.]�|ݽ�=����K���>�����/������gfwz9���s�������zk��{�7d���WC�����<�E�t��o��)B{O��x�'�>�����QJ�%	���8_Z�_E���=����}�<�����
^�?������7�O������N>����x�#;a�~��ۏ��:Z\p��W����vws�8�qӧ^ΝqK�W;�8{5ǫ^��!撎���Q��j���6�k	�2Mb�*ئj�L5&XM11ML�V�,SU�d�1j�L4LY&V��Uhb��&jM�-Q��1jMVI��d��Ʃ�,ecU�Z�X��&4��cQc�V�1�Ʃ���&5X�ƣZ�Ʀ4c2��Ɠ��Ɔ4��ƣ�bcI�`�&4��cY,bcLhcC1�cU�SYŌ�ƌd�Lb��ƣ5�cE�,jXұ��F5L`�,j��1�ƫX���h��cE�SX��Ɔ4�i1��#&1X�X�kP�U��5,ecS�ec%�Ldk+���,icU�,ic45�ƌacK5X��LhƦ5XŬ�ɌLj�jX��ec%����&21��cR���[)�&1X�c)�S��c%�-i4�cJƋLb���U�U���CF4Ld���K��F4d�F�,d��cQcTc��0��cSŌ1�2cbf�4���jƘ�2cb�5Zi�i���4Ʊ�6�b6b�ڛG[*){� ����+�N\�����;5���|�O�~�W�UA;x��.\Z&��ǩ��=g_̸�x��Xo>��mƼn���od蹎�j�?��ǋph�''�8>S��������{O^c��]S�|�ǫ�<����5��q�^�6�����vy_7�n��Bxz�R�|O����O[����ۻ�:-w�TTN{�{�P���>�j��/�~[��o#��}%�R��M���]�^��>���	ӣ�x8[Zs��UT'q�.r�>ˀ����oW+��Ÿ�_s����\���;'�73���,���P���]^�����4o?g�JܹW���z#�휸���W�x������Z�R毟��{�7��}���Լ��#���/�v���P��/�f��?�%	�]
^ދ��{<���?5ι�����|.#��Ź;n��z�ח����/)��;}�O7.W�ò%	��<N��=np���l�./M�r����؃��>-ӓ�p��|�gJ<���KJP�r�|���]��YK�t�^�d�v��<�����������u������u?����2�l�:x�������)�R箘