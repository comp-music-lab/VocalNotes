BZh91AY&SY�[��\._�py���������� � � X ``ҟ��        @  (  v�     � �� h( 
{�     @� �(�@g�  (��=!��ۑ!�دM	�^*������|�s�����x)����s������u籹��C1��� `Qa��IɺΛ�k�x{r�����^�0!���*� }��}��=:4zȉO�]�ͦO��v�zz 8   0�zd�%H$8u�Jh�wqӧ'�D�@!�E�뜽�䗡�,]���$�x��x  h{�)�Im�dÇ9��(�lLf����
H���5�<7N:s�h��î:rt�'��:�M�@��=x�PSٍ���d)Tn䊸�#`k["F��HP���e	
|> (*        �� T�M i� ���F�  dO�Ĕ�R4a	��i�ѓL�M��D�2�T�        S�(URA� L�� a���	=R��S@��CC@�d2d��U4�&���4d��ԏI�����L���z�����_��ɣ�R?�|Ȣ"����*"�j��!H "����}��>'����]2DP E#Q?��*�)�`SlD���)�"�J���~�l�>����מ��s�֕��M�S��;�@ �TdD�e<�~b�e�S>�ϳ��ϾŜGv��(�ҟJ���,�ь(Ԣ�<��_������'�0vÙ�Ǘ��I<���7�j�s�+Q�ݕk�$���gB��0��I��@q7/-o>"Q�F`:yx�Dp�����/���iۧL|;w�S�+�eנE�N��7\}�̛��r/�8��{����ѯF�W��U�� �M� ��zj��~�X=�b��߃8�o�+%Fգ��n��1�oi�b����F�Ӕs�l#�d��PQ򏓊��Q�-yFH6P���\t�Θ���7�Z5�k�9�6�Z�E�Mݔ`�K�"�t8�Z!�.�,c���-͆p�����G��7�b�DOui�a|�{O1ו��qQ]��%�-�l"������o���K'M	��K˓:-�B���̶p:���D�2��ۣ�f�o��m�ҵ9��l���sf��Ν�7\k��9��.L�`��JboqXtY�9�tb�t�������ݝ`��c�9EPez�S�8��H˘ɜ�\!V�ֽ�=ג�,���mr�aǼ1�� �8����Y���v�wVIU	p0G���ǨvIR�^�`;(�����׮q�b�$��fՎ)�Ӏz�-cFs��}'�-���ή��4Dg$p�v��v�u^��4� q��v��-��98����q�OYx�b�.�Tf�휉��뇭|
:3v[1B0�g�Hp�U孵�=G��B��tޫs�䞁�i�n�ݷ�x�.��7� ^�%Ē<ݝع��;���3^;W&����m�g���|5#� �i+���V{��~��5f�{AjK{^9t���s��̵4�s֤ݎ�v�t��⛝��ɰ�ð���ĖżL|yl��F;�f�(bd	��R&���xt�� {uqk4���h����i,W�.��E�EJ��.u.��t�S�;����mvŚmä�;3�-1>��Ŗ��i�;)Ҳ4�vC$�+�`8
q�^P��s���:�N�j��n.�G�Q��:#�Ua;ׂc�Ɔ�$��ٹ;T�z�!�.\���=��Ȧ�BೲX83��C���C�����x�sт9�u%��Z11y%u���X�7Dٜ�o�uzS;؆��Hw�;�8�+���#��/+1vd�z����{!�"�$��Z�!ZxI����,uoB�zw:���ܶ}������RQǱ�԰T���p�צkf���]�{6�1����z~�Æ��%�"N=�'��9�p�'���3cj^l"&���;rS��X���[1�-W�1,T�Ӽ���I����O-���%IU��×�Loi�qk�ǔ{ko5��ó�a�;79hz	�f�i-Z�M=������1'zo<�-YkM7�h�9er��n
��L;����Q��N��0��G��������O@����J�Rc�v+��;�f�����gNT(Cw�G��K٧�k��\р�1�r+��+�׀pu���ph ��/�c�c�	�i ��Nz"�8\6;��+��j��S*p�}Vjy�0Y\�7]�-����ͭ�M�ov��.���^���N{iǋ��;{�sxnk�$�[{7Rz`[gPd�z����&!�v�ri\Y�t=���r����(��w!b�����I��xj����M�ۼX�nڼ�4r+�L�n�Ӊ����e�m, ��Vt��eH�˻���Ӛ�#����wo9�7lI��'�{N�s�v�GpG.��"�{w`�ᑶ(4�������㫁ۍ�n�Q���-�s�<qCC4�P�ʞ;he=ۘ1��b�Ǹ<Z�[���j�}�1xw:�^� �75�-ɺ�]���,�}�)�û��2�>ADG&�׋�\�S;z1ZP�
�ٻ;K�A��9�G|;d���Zn�US��g)��� 7to#.�,�yQS�!k;��� Yah�v�\o-a�lH
�yGr])e����ۜ5�朗�X�)q�J�����wBfаK�wv乨n]�.��yY�"�q��"\��vׁ$;���G��ܽ�g{S@6Y5�c�Mw-��R#�;A��h׆v�G=�>�C��+�#۔�"��;R�F��'LJ����jST��CbY�ɛU��J�8v�.`q���v��/%�[�����G!�����V2��+�kz�y�
�3�rWrmV��\�`L%�9��7yE����R��U��Y�_�gf�H��ܓH1Ǹ��Y5��%qŃ5n������P3R�$��gS�Ź��v���J�AٺV�z�;>齈��i���<b瓯M�;�Ã;��vMr������j�]����f�т�WN[�RB?�컚�n9�S*� ބy�j^��H��ۻ��=��^��p���Wos�	��B������7����=��̆G������vsP6P!��5�^��mbh=ș��Rs쵳�:!,n��tt�i ��G^;��g[�͇ٸz�{v�N�7�S��tӂoN:r���H n�h�o���Rm����a&p�up�t��S�2�~���Ex:�l�pJ6v��4�8E�.m�3nݸ1���i')ӊ%ڢίz|��J���{�|Keό�V,�N�����>evڰ�nnPݬ �� Ȕд�k�^3��=�����z��~��0�χ~���~^>���Z2c��_�W�W�1�]g,��D�n	�� g��q��#����<'k�x=t�7[��u�݉	��#)t���im`9��s��Ζ:�;Pu=����&��b��z9�Q�{n[cB���u�������**� D��X�d�:%튺���ˤ3�rEs���b{v����L��g�˺��;u�y8l�f�5��b���֛E�s�s�����ɓ�Q;�ɠu�r���)��s�n�d벋�=�S���iT�N7f�]��tC8��Ɲo�0�`�2���J���T�j��+�W9w~v>���cq>�wvJ�fTh�@�>^۝!��z2��d۷��h�s����q��8��'-�[��9�Yv�15Uk��"Ŋ��ۆ�#�t��\S���9��Տ�}��lu�=���g��kt��t�tQ�y��!�����1ø���jv�;�a}�]��!9�mtn�he:݌.x=��uZ����n�n���rV����Lf�J{��\q����� ����p����B�=�5�y�y�:���ѕ�koZk��,��vs�E�]�Qϵ�`���[uWngq̜�Iq]���Om=�:ѭr�]��uѢ����S��9�m����{]�c���z������Qt�AÓd�ծE��vK�-�[g��Gk�;sE�j1�q�絫�l�	� C�5�<Y�-.۷�z�h���9�؉x��qm��I]G[twMOk���;l��㷞����ǎ�+����d�Ґ>�L���:�~q��v�F�K�v4�óu�^ОA���B�8�xZwQ��笚Q̓s]������m�)��B�P�����5�"֚'c��:�qs�l�>�뇭4�m�L��X���voZD�{�7m�5/`�vշfu�I4h�9�;�kEqi�3�ֱ���G��;jM�ok� �Wa�wf�ۗ�ǋm����;M���]�w6�2"�p��k���^m��Aۏ]v�!�j�����nlI��aݶ�/����.+�8���v����9���q����)��q<-���v��i�W��E�u/Q�<����=�.[���=��}���l�0�R�T1�\r�Ui#���3�q��l��� G�����ي7Y���R����ཙ24��摂Ԗ,@��>2�>z��1�"�l�-N�v�S���Gj5���x�������6ɯa�n�	\���I�v:��SOGT�n6=�ƞےhn�6��.�� �t�-�Jܡ�\=8[���ݓ���4�t�s�0��M�Z���Y�Hu�<<~G__n�"���k5�OYԚ<�җ-Ϋv�o<`����n���%�
��;�f[k���&��8D}�m�ɹ��8'��hu�hvEB�C*�S)����7jw�;gnb^��Żp�n��h9�o���I��Dn:��4�[���E��ӕ�lt��Ț"���n�w}|��E�΅n����s����-�%Tn8�q����	F�g��Ys��\:]��N���ô��
�vf�C�kB�����V0�I�q�y=o���ܼ����C�<nP�c��v��Wa�㞋KQ��l/Sa�N��VZ`��;N�A��=��]^TQ���m�RUn��'���מF��W]��<nh������m�������v�y9s�ew4ܧN�%��!t��z{U�N��gr�m������k4n��H�ǉ8�a鍍m�fr'��u`��g[�5��\�����-8d�iЊ�0͙�S!"d�p�a�[n�Zv�5��9�>1Znu��x�,��/G�����$\.7j2R�g!t�s�c��+��f�.8눸H{N��O(�nb񋗂�%^	W��\��Q0��ARg��k"!�~r<��?����/���`�7��_��Y�WmQ"��4�6��{'З�pe�%Ռ8U)����=]��}}õl�Z�<�t�]Ȃ���]ٯ���Pvd
�_d�����-;C*?xɗV!���>����o%L�t�n]���w�W���;��ʾ�j�B�/=i��o{�|�^Q珆jm�yϑ�j�Sv,쌞��q���< �
S�}�F۪/N���;+>�����ɢ� ��)�\i�~�:�����<�Ƚφ���X6<T��'�;�N�j�o�3�GӞM��y<*в�ך�=����aX�L�ʲv��aR+=���=<���ǅ@i�O�v�}��uMݛ&w�!z�`��q=��e��}5H7���I#�Dw��}���v��z����7ܴN���$E�v�ދ�^��o�T{�:������y��y��kp���ms��R�x@}�[K����3���uN6��p�L�Ŭ	�x���1g��Sw5y
��EȐ�(����E��Ї�=]w�f�G��=�l��郼�Ɲ=�oq�{*0�^�঴�`@S�;T=DM%��rf�{9�����e��wS�!�Q������@9_@���w{/^,���H�xI�N��C�<-�����|����]�c�zl�m;��d܈��f��:�בz����d���6�.C�"�{�}2�5��%&k�r��4�n�x�*�rr���Cg�9��w�G2m���� ��n��1���<���ޭ���z���נ�B��|�
���x�筊�,<�:vs�U$S�'�D�$��v�I~!vrc�v§�z���\�_Ix��ۑ���pѵ�t=rc{���@�����ҴS@fNys�o�њ�9�i��+��Vw��;�3y�=n(xMM`Ry�h�yI�L�S͡����C�e~�����k� ~��f�/:8��+l��=���?DLH��{�D�~\� ��/C�A�Ǫ7J��m�}]{0�j�cC^�0��m_+���_{�W{%�[�!.5���;z�����qҼ����������&ˡ�+�7�=>�h���KV�.=�0j7�90'9e���-4�n������}�k��o�I�šn1NO8.���Lr�'����w�Kb>]�>cN��r_z��[�%e��Ou�>(�z��`���L� ��/�9����##aN�엛d�եC]��%�Jī���W�k��P�MmJ���(�M���R�2�1b<��W������^�ݘ��h��=���euKa��x>e������پ;Q���^ѳ.^�b������{�K��y�(�C=4Nɷ�i��
`^�r��q��g�2�Y��o�����s;�DΏg�S�
s��lh��w�p�fn�S���-��=7�{��_�r�;N[���4�Ւp��m�{T*b���>�vze�x�-��B4=�'i8��1��^�d��}����;�M/���Ñ{��[�L��7��˚r��b�K9��3ĩ��n���Q�]`l��9�`sSy1����9j���gHj؊{-���ξ�)�7!�tL��=��6��F�]��v��5���K>�l�gd�z�����F�k�ay[t� o6��|O�+����T�,]�G��*�����F˿,��ۈXF�l`����g#�𫼷��n!ӲVם��ե�V�R����y��/j{v=�I�������c1�r�����z�_s�X5q�ݞ�}��`� �ݵ�l���y�r{�R=[�3�ݽ7<r������c7 ��-�v�o��{t=����Wc\���F��f�;͇ϗS�����:/v!�=�sy>���G�?b�u���Ӏ�SA=� �0����d�)����v�q�[�wVG8h�2�����k��Q��op�
�z�|��'�lX��{k˜�<��.�;s��<�K������%&��<�藪� '�#U� �+9,���$6�׳Ϝ����w�ʔO/�DM���e3�"k�2�b��B�*t�l=x{��f
���>+�C)�>+6�nn�9��N�YD�^��^�+|ߏ�o2���;���
�e>����·��ӛ��Y۞��f�{����MƏ�C9J�ee���w}��V��*����\�;���0�e�=����-FܓC7����G�k�b��Ժ�7��Ѿ�l��^C�*X�h%>n�f���m��卑���	�|�����}���f�V����d����Ȃ*�*��C*YY�+3 bW �|�Q����Vyj�� �q���iվ�˾>N���ۗ�w]o���w'��v�=-��ʁ��Dk���Y�q�-c����'˾���=�83�����i��x�n'�)=n�`b�ps����
���)�t��ƧpZέ��ɼl��*�hVc�X-��iW��A��R瞸��_a�������x'���6���>�dе�����<�7{�.q�v$��,��4�f�|1&y�{4�����s��<�L�u���)���N�������[�-�U9��ծ��s���L�њPέx������u�>U�Փݯ��g¯gwA��`"x�o���3�q���g�}`��}_��$ Ha?ߏ��8�� x��`y����%׎1sK���Z�i�V�r���!��P�neU���uܚc]���;LC�G#Og��ZG�Y�Ż�#�����β��{q6��I�]3v����Y�g���;����-�%�۫����Ӵ\�tY�]��	��WIۭ���^���vaq���6��f��N�sϖ�.�Ӷ����v��3A�g�;A�cn����z{�:��q�Dp�\p�#�e��y��˂���[��c�c[n�NN�������ڲ\ㅭq��֭�q�F���=���u���r=^mt��rv�qs�Ϙ+��
�Q:z:��p��vK\[����8�Ǎ�(V�=9;�1��:�m��wa��0dw��uu���˞8�Q�s�)c�5��]O�R���sZ4i:M�������sӼǇ�{��V����W4Ϳ{�N�ӚӼS�ܙ �y+CO��t����$WV�Z��kLܪ�FWk@�����=᛻��xr��w4�l�n�v]mch]�@��^��1_�����m�k�Rd᝽��m�6������UJ�����b��_tzH߉�f�5���8,t��|�y7�\��Ͼϥ���O��]�v��
�3uk/m�_�&�O��9$��N�����ϓА�6�cO4_}�V �}g����^�ۧ�&m{u\ݛ�n��p5��֝a��\����b��m���\l�ڛv��ng�.2�p�.ɮ
��^� 8�>�=}��ogx5$oI�9���5��1��g?�К��cy���.��,��]jM�G��h�d&tʼ�tǼl�B��y�Na,�w"�M��}�� ���x��*i�u�A8�����X��=}>eJ5��c���vv�����^��෍�x�j�����ǅA �A�$��A�C���Ϋލk�4lbɞ�#�t�"�<�	��9������V�=!��γh�z6��K�HN�%3ÿor�H��p�Y�ګ�Mh,Ӎ�	4}g�@c����a�R�5Mǹ�"s/�
�b�q3�K���W�=��{q����]A��m�nK��1��O��6�u'uޥy_p����,�)���� jT�e�"T�_l�/�INd[��q�3���TFL�x����j�.� wT��vgu 8C�lH���ҥ�����j��xϊ�Y�v���G�$�AX�S�I�As��awSj��]� 	�äu���i�QK�([[z�K����/>�.W�#55G��ζ���&l�gF�[����OaH4mbɞMzP�1��á�V�h5:��R�{��R�ϏDm��Z"srI�>E�O���m��:>5�<dy�m�q���\\�x�i<��C-��|7��v����nغ��n�tI��;v.^Z��75��S����q��ﯾs"�䭄RIQ[��Q��Fh��4s��6���{S�3j�&a��׵�
"C��+ެh��>�`�1~��𑐄�΀$:p]�;q6���(BU*��u6��W�ZD�7�V�<n�t�49�m�W �Bl����ގ����1\u�9; H	��#8��W�n7-�3��,�x�	�K6�	5xV�B��!<�۳;���_��g�����/����8U*+m;q��gp�t�n�:��8qdhٻrLNg�E��/(s�N����U5F�DS�Ӧ"^��L����.6�7KV`p�F�I$� �J�V^��_�.�Y�)��jkr�x�g0�f~9E�%���qK"���,NH0�
�'\�\yP�����
������U�a��x����ef�:D�3�[r�%-^��Pu�fNݜ����mEfC��E��\�nSY�c�8�; �2,PQK�ץ�||>���>�ܖw>Ȼ�x��ƝSv�ZV�5e#p�$���� g��T�X�h�Xڃl��m	ΒG�i�P�k\ պ��9��N����%�C�Ӫ�P�u9���&ѧ���V3����h!���ޭ}��^�v9� Սn8�ʤ�ۂ��p��v����^lT������ٍ`�q3n�\r�n��.������@�#n���L����Zi��I�6Î<pqۺ��6��&�b��4��a-��}�ֳ�{�L�_r��Y�!��]Q�#�F�[�b�T+��^ �rYӖ��Dd)��Ӫp��Eŋ���g	k����,��D������ֻ�/��)̋���#�����Ċ�d~���ܤ�4W��o��^�/^|}��!�0��y��1^�9'$��g�i�x����#L�@b�&V��Cmڧb̆��B�Vl�?qm���	�*�#�b"�USx���:aֺ��0��E�U�!Q*��>ڔ�����\��l8�}<1��n�����+1�Gs���ќ5ʢ6���&�x�`=5/yU�g��<��s8.���A7ٗO���x<�C�� ӝ�/	��� ���n��;5 ��xP҉�֥�ʝ�ջ��]}}�_
�D��^��y�O{1�9�Gܯ���d�x��f�0{������8�ޕ��t�׌t~{�C�N��GZ}�ݜv<@�8Wʲsq_U ��
�	�^՛.{��H��nub6�K����ë�,L��L�o�x��g�exK\�#t�1�߽堿3��5�8�TV�	�;9���T;��qٍ��33[�Q�[�T�8�d&jN���B���K'�͈6D{'	�q&����D�S<p ďA�f5�P��6*��qmyf�t��=�hՃ8�\x���|���bˏT����S���Y��
�۝̡28�s3�$�W�2��ss[;[�7�)Q��{�W�zr������W�D���(��C.9h�h7$�Ԯ��D�<�@o=£3�3���7�W���xڎsݹ�e�8�t` e�/�px�}[���C0��;�D	�JA�}oV��*����i^����=
�]RQ*�i����0�q���ĬȮ�=$�.�݋�)^T�͡���v�0U�ƈ�Tr`�W��)�)�� 9���UWuyG����4�t�Y��b�$��^E��t�w�Z�����L��E�^�C��C�BD��L���l�ɑZ9��L޵�賦f�I$��	'���6Q&CK�ޚ�������yz�z��w{�,N�%�%��O�|R[S�2K)"�K�L��XX����+\A�/x�z&	yS��tLsH�y�u��V�ٽJ�^
��
�r�r��!�����g�J��`i o�q狵$]���Ѻ�����nZ�w8�&"�K�w�7�pE=�Բ+q򮧞�ڪ)���3;A�oZRw����>�YU�ˉ�6�ó�>��ίN���u^1֎�]����ݶ�Wj͇��<�27ۚ����&�)�ٮ8��k�;����ih<\�x�����O�q� 7�]O��ۛ�!ˆ�	c��0�X��CX�`i)�\S��Z�;�kd��Aީ�1K�i����W�<�nԛ㚙L�9�@q\K^BC]��).}s�^�b�^ �17�-I��"�7þ
�*VT�kt���k�L����.�La6�����v#��a�Jj]�1SĮ�!�������坁�k�B��\�^�JɈ�M�F\?=̌���q�W4����$��WG"�b��-$/�A �I ��Y)�BbR�����ѷ�9���������E;��&y���.����M���WYC�ot���%@.5���-I����$�C�;���"��8�o��$N��.��>�g��DV�%*rHX��C����3x�L� Ƣ��%�!���b������q���ţ��.Г)>P�Sy۝��$:�px�%�����ʓ�!;k���MeF�H1Y�p��e�b�DRH$A$	,�"�"D�d����C]�!��2�^�Hg�)CWX�u�bp�Z���.jM�֥e3 ٪�t�bԐ��K��S���w��@��:�1	SOX���Gjf�su�hHg�B��0�qM�;�5�7.�"H�tv1x�IU�Ա��P��s[%�P��T��\M0W��=�J�ԛ㚘�b�xD{���^�kq�.�5A�>�ʻ���A�j��,T�A�$H$�O���"J��EQ�!	����W8��̋�tk8�+��Is+��(ٌb�T��mNU�z�0#*�e��|(�z��K�����U��+�t���v����X�c\�of+(�x�qT��Q����RH5��UwW���"��,Iy�.&"TN k��;6K��]���st��4�SUԵ$?T��`�ǚ�(:�s�-9�Z�z��}�3�,⬮<�m*�e�>�kַ�w���r�װ���I�[��}��B>��K���o�똶;]f�Y�6��v�F�d��n
�m�ti��x���A(���4Ǹ���/�uج[����Y�������I�7q*�i��ꍌ�k�B���G[�V%�$|�s� ���Z��H\D�"�pnn��L�A�T�P�b������M�7���Ls(i N��.bTy���Ғ7̮��f�E��S�ӈ��r������2�5��qF��������a,b��Y3+)�����{����!�K����f�I��q`:s�)5&�nZ#io66�R6�Ah��SZ�qH7ߏ����ʁ5�4�e#M��F�H\Ĩ9�� +�S�]�I�$;�q3T�i���ӈ�UԵ$4q��d�2�% ��pR��Ò��@�1��k�qL�|1����g�w��El�j�'#dRKh����3&l,{ׁ���S`�N�wz9*�US3�� �s[�ݥ>>������s2yyS�Di�\����W:pS�1�Z�n�ͅ=��$�|����c!�>���,$Z ��4x�[�$Njj /xk7ȳ&��Ŏ�!�E��k��=�P��*��lN��^����GcI��H�{8X�����{�].Hմ��90v��9alШ��x-H�UǖP�����3A;��;��l˻�G:Rɨ���!�H~�����׏��xd�`����H%W��ǯ�>�/?���=>�1a^�W�u�OX�u�m��d�	�Z�zIEc2��^�5b�����G��ߑݰ�Ѽ(�[���>�X�y�)R8�3����rK%�v�1@��-�c(-vi�xcacb����d��{�˒&�1�J�o��|j�+vb��ht�d�͵��2�|�c͌S
�*#3�I��,�}�P�n��X��~�C}��+��3�ƾ��#
�1�������F{TֺOz�,W|�^������;"�u�����y�W�����x��H�瘓�j	@4޽�D|���h�����?qy�ߟ�{C��@�}��~�.=
�ԇH��>�a�`�]�x�ߌ����u��.W��2yq���}�i ��G��*K5�_���B���� ���\B��ؼ(�/]C����x3퇕��]��X6��O�2h���k]:�]�X��D{��Ncӓ�4b{2�{�2���|�������J����z�;Wx��#nbF�Z�-H֒��TL~&r���
�.ܡ�G��k)�	�/k/�b��lmە����\3�.Ny$8|�C�i.��;n�5��[��٫Il�oXMw�o���ۚ��B�-f���q�o3��U�$��3k'I�+��Ħ;B��N5��^#��lOb�lÂ�.�;<�۱a��q�T�nrg\���m�����r����::�hث������E���ۮ��]�-y�VH�屮wvo,f��93l���R4�"[e��R�>_��>ָ�m�\��ڱϝ˰��`�Ɯ��XG6�g�J��4�Q�/���PdLh꧟m㓋�S>�U��7f2i�d\�ݷ<c���P��v�÷c��JiÚ��cc��0��T!��ԭ=c�+孽v}�M`� bm?�� ��*f�'Z*S�����h��7ܯq�~�wO<�v9"ɲ �Z���:�Bf��vtX��N�4��n��N�����B���7��mf�Y���i��=�y��4{�.㚼6����an"a���ib1]+ܚ�O2PӡYU��T�wˤ+�u�.=���c`�H��J/��Z����;�)�tfӳ�8V��LKnP�I��Ɉ��{@�Omқ]�3#��s�X(:�����̘�M�϶l]9�2�7#�;����̙���ݎQ�۷U�Doٯ}�q���5N�G���d���Dqv���
ؓ$�M��x�����R�)"���ظ�����E�n3B����� ğ���;'<�����~�4�0������_����{YZG���)������
��&�y���wze�~�'����H�#I{��NE 㩢�9qe�Cv�5�%R��Y�T���R8 >��QG��	�[��u2!�7ZN��b�я.�"�3>>�<w׷������μ,�ɀ����V1�%�Z���ߏ������ ����̒RT<|<23LĹ��t�_�}�{m�ͦ:� �|�'^�a[+���5�cOٝp%�0v��::N?{��u�Xw��ټK�˾g�&r�q(�����1�C�{���x,�IJM���\Ҷ{�s�CJ8�<�`�-�];�Rd� z��||�y���0�M�$�� ԃriґ��F����D� <Ǻ�4`���� z�-�l:��^���v�9�EUDrKTRVT��U2b�L��d�U��뛹�f���3�o���\j�n�Y���77��
޵�ws�<a,W��5�,�@1^{�*�c	73[�_5�k�C;ь����
%9	���F0ج�|H"KA�01���{����'3&�\ >��l�ib�����Q*\�T Zۑ��5n5����.Uf��bOso�G���PQS\�2�:���QJ�s5\��p �vl������(а��T�:;��fs�����������;�Μ���=�j#eC��wgpkigg[L�}$]���V��6]���s��o2D�1�B��TMo��r�{k��E��<U��B���mX�S�0G�`z6�u�u�4b;7@�yB�g)uZP?��J ��ׯ^_�|yN�ǎP��	3����a8�2ߴ�y��0��F�0��	�۬#��K����ä�� �
\3W�}�5���fto�s�<Xi%���������]��жi�Z���z��K� �=i�i)+T��br6Z���4=c	I���e��c(.|���XXح�x4ɬ7UQ�K���5�f�%Hkna<��F7ctE�+����x����}�!�� ������;��H)��&����;�̛s�O>C�|~���\I�$��]��\):�.�F�cU3;��,PV̜�`_/��[m�b5�PN���ڗ�&j�t�;~�<y��q��Y�]��:� xz�ܘ쀽��W#��g��%�gw�2����T�tFL�W���iUp�D�צ���s�6�������2���1�w� cIk�l	C���Dv�2��w��W�;7��}<N���q�c]��k�m��6[1-����\���hWZs$>��������d�N��F�Ưp��;�3Ԙ*���ҫ��Pټ�躼�ҫ�9�nnNU��C�(_*p�+ յ�rB�yw�g;?�}�ￍ�04I��Z��($Ղ�?J�{���Z}>�g�������i�;�����ؠ�Bj��<&� 6B��l��wo�j���u:��*�k��Se^u1uʩ��6cYz�.;�X���o&�}U����<음V�p<c���b[j9sgl�<6��N���k�8��s;��ۚ�v|��7�|��[1�v�/`�W�	v뷎���Sְ�Ok�[c���w\�2(n���J����l�c[�t��FgO5�����{���{� �~��y�NuzXM���O�{�7���vH����o�`���1�����ɵ�7�7ܸ�1�^>�sE?f��j�k�^�#���	��*fǁ�73l�ґ�۵N���POrc��>��'�����  ��t���QP���g�0��6�S6�h�Y����a���b�*Ż�;����̅Yl�a��!��t�U�O*/|I,F2 c��˜��chQgs���gy�նx�̠����\&1`<���$�� f;v͡��M����l��~��[�5�Ȯ,c��I	,oIZ�\ʅ��kg�}����₱�4�,-��4�a&Ɛ�����H`��c��\�-��`�h�XOy��}��uT���awf{a�q�}(�=}���C�~؄�oȪ冯x\��+��dG����]����|`�H,�/v�N����`i�Op"��ON��7d�d�=�x�����{������w@���y-��w�sݧ'�υMd��þaw�漊�A�JN �vr;s��[с,Q�k�h�rV�>�Ce����ת�]�&����iǗ�Qa�T �0�ӫu_�]d�mW�.٣��ݧv���yG��|�u�{E�
%��`��@�����5���8�7���.72�Bhh�31.��M��Mt6Lem����`����Y�N���x�1��0�=��#Ĕ���ٚ�N{�E�� ��p�<��<�O@.=��`=����W]�{P.k��N�/���۸�/Xy%�߷52�<3�	�C���~�sϗ��q��H�Y�w���u|��d��x��� ���ұ�
�m�?pdi�������w"t�ޣ\��_�]�8^��2���>q�7.��vv�E{�{�FF�9��ޝ�n���}J0�qf☧����>�h������z��r,b�4g�|�����F92N��=��z�<�o3W�G
6��4g���a�jqǯ�t5��5����+I�X���q�\iaf��aT޾�����ǟ��-���Rk
�j4k6K5{�����HL�AK�_���73l��J~��}�V�]�Kw=+�e�w&��F���Nڅ5��V��TFLR���|64Q�1�[������>]3��zm9��ل�7����NIcs��.�+��߇���qr�;���1Ew�!j�$��\����tL�q����3o3T| �ؚ��#m4S_��/щ޷��<�{�j��P
8�%�h�C {��՘�On�N)����7aDfQ��7)��D�-��.tFY��}��3�~C�D��"���{`��gO����sɻN��D�������6�"��q��ösV6`�Vul��&�&��������=��v�~l���Av6�t��{��xf���'��nߞx	�&�-��O`��&�A�G�� =qAP��+��V �	�?ZR�2� {��D�u#��y��кR�| y]+�Y���ʓ��ZV���"����u7�	�u���9�Ѐ�7N�I�L�0k�*»G;����*��6��^�u����G=w��`��LBF@�$'��l��g����咃z�j� �v�f/�\�9����w)���)�E7,�� �tớ��U�I�'l,+T�
5���G�-��B�� o��]p8����� ��Z���\$U�@�I��*��U3��CF�c�B��7o6�4�OV����b6��[���=w������<}��
��j /{�˳�ߔ�\����㍧�ɕ����vZR����,��T��+�9n�<�zG���A��V́�d��^F%��1�@��6�pfx�f�f���A�₁�4�{��[��c��K-ao�2�}N:kf��9q�<.6�i=	�CHi$�	&Ʊ�Ys�pʁ��,5�?zN�q�	{�o�v(ړF����1��^�f&����0�����B���q͞��E��1��=���J=kݑ��OJ6�;#K�^'b�~ �x+�cis�H{��^d�o�x
�mA�c�ٳ��N�9 ��l�hV��VAg��޶�̷�m��� �.G�+�q���p����p箹������t��*]N-5&�FR�R��,	1�<�q���;]���؁*���I�NԨ2�J� ���o�\���1�@��~�{�����r�)�R8��>�bAo��t�:��EZή�u]b�
�E�fn�C�/{��Ԃ=��f@���C�k+�mK��֪�9���n�����"�ʙ��j�X[�'�3��bp���ȤD��8���!r��|@�0����I����t!���OV�R��CUӛ�w�mk���y���u���4�YFA�I��p����١*�� ,4͡�d��kz�q���~�[ԡƇ� �_�����1�-���~�^�č;Y�Q���.�3��L�#��#{��4�.�ef{�L-� x����҈��J���u�)�'�U��6hѰ�S�$k����؊ѹ&���~;��ntjx Fb�̣�#�S3A싸�|��N���_{]���'#T��x��Ct��X��~�X����lF��n ���y�ݼ�;Gb�V��ہ��%�P�jD�L�H�L�]��U:Gx+���#����S+�~��b��%I���\θܓs����ۋ���3'y���n�c�#��	�9t�"�����/[��;�㓠��`��6�,��{�yf;%:�3��X!ɌK_��;e3T͡�4�p�u�<#8����7��$�פ�9�Os10Wx�V&C����۾ʁ�4m�+TF��ǇܽژF�wp��
�}�����K|�8�鎺����ǀ��a��.3ea*�ʥ����c��5�5ê`lD6�<E$�g.�."����4����O�kƶ7	�pe��g�������^��(j��[Y�]9�%;�����XSK�z/w?xpө�Y��>����,{
D����o�g"Bĺg�:^|{k����n��_�����7!ܞ�]�����[����<:o������/�����k�bכּ!�&Jɣ5͝�����������~���u���6�1η�=x��S
�[���;۳��Y���md8�Ļ���;I;S�2])D#ٸr��c��+*�=l�t�๶g����l]���=��[��h�Zgn�G���9�q�ѣ�LPիݮ��^k��G)�>��x�8�rj�(�%�{���-�9��qvnu 	�v��c=q�n�:ݭ�[��H��k{{ �6z=���\���R�t�E�`�)��c:{X׀�|�����v��b��`v6oJ�mU֙�*,À,�]���mv�K� pI�b��e�V��R*dl�7c�6y[FK3����`q��Od�$��秴WN��<�ź��8� ƓBn�� ��k]��μZA?A7r��rh@dh��q�b+~c_��m}I(�āa�)�����AN��{��p�+��#��������>�F�b��ʒ.z`���g?jl��s�d�N�㫷O�(�@nin�eu{}������N���{�L9f\x���م !��4�߇����z����e
��g��(��LGj��7~�y��>���˚Wi�wl}�ŋC���l]<P9wV�i�Z�������D�ɼ�W	ڹ��e�HŢ��7Z�䱋���ۜ��e�eB���.�b���"X;O[��IB�G�cx�$�ȝ1*k/LhM&��o���M4�Q�KR�42�eJ�Ɉ��Ӕ%��f���눝f�ҳ�^;�?>�|j��ch�UXC+��U�s$�]#������f8����b��w�~f��x��Xn`�kݑ�������5�k�o�RQ47QpH�S�Wlo	�Id�O���R_w���L_m�1$�p�%�7��r�bX]����q-�׆��]�P��z�|�|\�̮iws]vn�;�"Cx�mA���IW/ʡX���w����~�cE����}k��6�x_cZ��.�x�죍Z��*������B��X����4���k�_+r�6��f��6֪�n.5mP!ȐZ��P	L�2����j��<��ވ�yϱm��yLxb�cHd.,T$���p �xM��K[��rem��O}�cޭ�Mˉ$�1�B�SZ�q9T��I�E��0���#�A`�Gy�����eZ�2PwY�0ly�������l ��C6�1���GLe�[��W*.�Ȧ#o+��`��FX!��e3kR%"�("HDQm�@�hv1)h.��G�o���)]�������ZՂ��U,���z��D����nH�}���K���S|o�'5$�L��9��c�)?yݢ�mv���r�8��:�M�㌟��HG�1V���ڇ����#�F¨�tIw�c��'gb����m�F��ӣq��{=���`�v��V���G+��=���r�D/k���N��<7W1�0t��>;�׋�;��-�
\�ãC�/,?����L�x �sh.�XJaaG`�ד�#9[�J:�B_�k�x��ʁ1�v;��b`��}w���`��c�M;��d�������>��8��+1ji�I%RM�jG溒�����ꑃ�Sl7<*j�빦�K���FĆ����1�����k%d��j>)y&��M���#y�`��b�}RjN�Zí�h�n�4�J/�w;%73HXX�I:L��m)ߩ��]���aG�&�P�΃�h�W;�f0Qna�:�f��&{��iM� h�s5�0�Z§'3����]�6�`ɖʰ��q�+��1q��-�&�cf�~a7#��[�
��aYy#�5�^X�ͅ�t�:cz����[_k�9ch�!qQ0�ݠ5+v.�Q����s/��f�Ѻ�x�������]����3L�g���k1!�9d�_�[�����֭���lȱ1Mb��[�4�G/��*F^];��AI��I �|v��ks3��tx�L��M%���A�Rp���r%Yp����>}#Τ��$�/�����o�L3(�4�ι��33ť0�^��BJ�(C	����D-�"�d�$3��"l�\M�=�D�1V��5�L��� ��}y�
�4�^���-m�ۮ�ɵ���^;p��b2yu���4�&����gu�f=%X9�U�V�=S��r'S��Zx�����#���v8��]u�d��i�j�9�Ek Z�+U�9d]�m9�Y�sft'�V 0FB�� �uA��h�� �m���,�k�-T�0C�����`S��)� $f��ߋ�H��G�x���[7��:�(Kb�.�2�ꢷ�nr����+���b��2��Riֱ��x�ڲM�<=����5�߯��)&�YP���wx�gtfl ���.J|�$Ur�,Te3X֢�i������jVYZ`��4T`�wv�^��ol�ƣ�}�n����$�iO��l�2ЪM��ٴ	��lvԪ�Π�3�qݍ�S=1,PPwU津jY?l�?�)t�]�3�6g뎞��������tĤ�f��p���zb�B��D�Qw�\5,g��͖�$v�uÃ/�߽����z�a��zwr�ћ!��$߃��ּ��������Z�2��o��]ðp���x�'�-f�9m�8JsM0un"JM��J�u91�5M	�B���,�u��ڻ^��/X-����ȑ-���yƈ9NmeB|z��7v�}9�w�������A׫����>螟ٶU�G�{}!������t�Ks4��H�hȜ/�Rq�Q�Ɲ��iA�j��ϴ�>��>)�Q2À������o�vQ�wa@稭f�΋�0$�N\e�!�ѥnѺNًՄHÔ;u�M�KsJ޴>��Ι)�Xt����T����,��tK��^��\����9�M�yR��b�ax=��^=b���t�O)p�ۺ3� z8D�Kf��a��1h0����1��C�?<�]S�'n�?���tp�G
-�̾+g 2�:���.e;��jf���!���}b�.�SU݊j8�;�qJ��4	�#��3#���ڄ��^��i"���yÈ���V5�_�'ړk���A\��	��
��4"�
���8^se�<O4���ꙹ"c�J�x�f0U���o�qPndfp{��B.�����<k*�v�c�`�R5��ZZɱ�Z6�^b���`�Đ|���$�H�"
D�H�\w�3[37l�<ӿS6KG����$�v����n��������go��#��Jԏ��g��f~�g���h!� n��9Q\��w�ʧ$��`��Y8M�Ƭ�;�yh�n�0��۶A�Jl��O8݃b��5�&����7v�b���bb�q5"�j� w�]��M���7��C�>�N[�m�ԁ��w��z��x�F��s���-�J<��b.��܊��s��k�e�y�;Ü��5ݫe�� �B~��!\-�[�n�u���?��kE��ȫ l�p�e����O��ä�a�	��ucz�棫y眣��TT������ �nA�¢k�3�}l��4�P4�L��9+�O=����P���Xc�|-��T�Yn&�e�8㺻""�r�q|�#�eg�H��SH�Q
�:[��c��	�Ǻ�̔v�y^;v]�r���db��ˡ�5�����c�Ht�jZ؆�Um��Y,���k'��)�={������3\3(�4�]t��.���R�}R+��*��6kbPn��H$5y�Se��������`��0с�ok߈�[��ʳZ�󏚑��l{i߲�Be�!�MЫ�
�������kh�\q�{spLP����i�n�����$FLx��lԔv��;��6:S=��լu)>3?p|%�1~[jit'
��c�ILu��ֱ�%F���w^�S.��n�f<�AF��hi	�@��&��i�	6</���[�;�+�_�}�=$�繦YW�J��du�2�]{�oR7�a*h/<��M2x�<��m��(� �'�1.k��s���8����o�w;\�t�W��LrYSpv1<͞
K�cx͵�o��֗Q�/3xU�	���V�v���M���IXgZ�LN��F
�GS��gj�8���i��֛]��90�,'A#�DK쑯2�.U�ԔT�T�%��2��G�M�����˧\蛹��z�_�nm��a�u[����^��us13i���L��hj\�٘��l�ԞԝԛH���+��M��rqaq��=r��.�`�{�b{�_���B�Jd�G�2 �3t3X�A$��rK���`
�;/h�w���`���w��v����2w�����3b��Y4�p��h�{��0=n&�/O:_o��cbm�@Ǆ `�!�6��<&�hcL<P���R��j�.��\�	X	���3t�s��3����&&
�y��;��dT�c��N�,�2=�����r�D䣄c �b%�����<��:y�h8�/�s�n��rbb@	���I`f�<Qhk��T�8�o1�KfЈƬxQ�m��޼�'
��;��H��\�8�%�x�S7C4�0(�x�!%r�	�z"w�f����Ҹ�6;}P�7�ݒH0f�m�F��m�%R�lc�Ӹ�;&}Ӌ���kݳ�zG��V!���#PGk1�k����	��\!��K
t����X[����i�yg�YD�R�5D4�9�/&��g��(�	H���ц�cl��B]=����t���+}���X����U8��&-DTm�
�7��;���%l%P9���̠�՞����l����vd��zzJ�=�[��m{={����0Q�f��+�n��wq3��}�q%��<����Q�����n%���|(9���YƢ��z�S�K ��yo��\}�`_��쮠�zT9Ӝ�R�E�WE��v&r3Zvŧ�S-�#��}@�CЂ��ⵙ�;��h��i��%R�t?����%��ՂK��Z����`��ˠ�6�N*�۠��W7�_�MC'{5���?W�RտV�q�]��{ӳK:�ty�|���N�R�j�l3U<5�	@B)<TK����V���j�vʱ�,�]�4�V]
0SFb�:�3N�rN,�k�6u�+�(��~�V��V<K��>�(؅�՗��j��]o]:,L�k�.��`��v���̅q��X�<�c��v��|\�=q��u���mƗ�ͭ=\�\����-m����jNѭa�mu�]���F�Ə	�Z�rv�bx�j��6]�5��8|����k�c>r��9�;���q�hm����mKҁ�h��5m�s$��PQt���u����V�v��ݻJw�56�n��q�-*";/l�v�<��KI�u����5��U�n0q�ܼ=���v�[=
�i�Ρ���8��=qcl.�ӊ�9�0v��y���m��7O]���\ݴ�=&�}���ƹz��f��k�n7��N�'��^1.υ�l�Zp�\��p��Ѹ8Ґ��s�*��s\�	������?q�?2
���E���Ǻ��&�V�s}�v���Y�V,Z�<Z���͙+��ۢ<��v����Gl��<͏ܽ3ݨܛ���PY�p���i��jh;�ES��Φ�a5c�jEz"xC�w@��iır������z�
(�ۘhǇ��WmŸr[:mGr�L)@Xs��}ڍw����5��c^�)�&��x���2fa��ڣ�0����W k_&�殛���dֳ�q8�O ���퉠M7��I�"���v�\�
��@gn�tRl�h}<{V�� ^J����s�9rh<��2n�m��wy��y��9\�]�N�����li0�h�.I2�-)S#��)$ER�ji�+\�h�'{�T!�7Ycs������G�q=)Xd�]���wSd�rzRX�o�ZX��J@ͱG�J	�Ls�Ig�c���盜�`�UdEm�ԭ��J��GRd��=�G-1�f��bu�r��p�s|�#K�K�����a��ɼ�Z9�����w]Φ��30cC04������M1����n*���&-g���O�լ�531��U���d���ܑ�b�<C)&��쌈?1Ϥ{���Ў�����CZƣ*���u��f���J�L�v�yQL�+ On�y�ԏ5@�4�����=I-��7i+j�aj���M��ne�*��V�h�4&�`M�@�.��d��;��_�>�xQF�Qfg*g|���.�iK51#��A�^�I=5<s����y��qA¢R�$Ptvѹ�KKkZ��H���z�%���H�קp�MnOs&�<��C�M7�MIď8�d~�P�< s5K1=ɣ����jl�oٛ�Fl]�{��������n}�ƨ�C&c��wN�R2��:��:䎥ӻ�\ߞ<;����������勫_�'����=���#N�"��eN��h㪆����Y=� �p�P'�&iw� �z�R��nr�i�X�s�݊G9e;M�Ч�ȇ4N��2��� N��C1�Ș�{Xk�ߥ��A�S� 7�˗�!V�@����1=tWn�a�]��:�`{Y:z��p�ti��"���k��h,�ۮr�S<7U#�7CĎ	N����<���\���i���9�ݺɉI��ؚ�:B5l���@�h%
?Uʹ���&��IB�G�z�VG,���؞���϶WS<�"��>��/�4����{�oL��%����5ř����;���NjcC�޻ivk���v��mcf�^�
U�3I:�6xW��*�s���f���J��a���]�]����W%�M���ޜ�ŷ�'��f�@�&�I �� �hci�F4<�����gǼL�Gk1�k��K1�}GTÚ�A�P������ê��Է�[����4����9���2(�*i��c�߄=fG���-�=����Or��FJt�� )�=�3T��jJ�r���+fv�7�b�6�5"�͕4L�IZ�r]=���hM���	N�v���J�w�~�����ǖ�,�8
f0Q�f�+�hk�&Ql�=�~+zd�}�-We����I$UAI\��[dc���{Ԟ��ԏ>��.��|���>�g
�׬�Ebυ0�@.n,L��ep�3k��c��-�n&M+v���m2�9u��&��t+!�d7�w�8ݢLN:9ܝ����nN�4��.�n��&h�n]��'��������Ϗ;/ǜ~Hӗ�>1�[�k�hZ�D�R� R�J�B+��{zMCo�b�Yӆ��&'�<ID?3��w�Ts���k1�G=�FJ|f~n��#��\�f��*�K��}d�yr򍕞�w<Qlf*�sf�p�;<���k���x�����]].j��B��T�	�\�[��E��;�՗�Mx{�������Lm�Nf��Ý��]q�eNֳ��W6x���Vti�K*��m:6$4 �7���:t�.�B�p�h�L&bFM1���LN+[Q�ԂB1��PI]MAUSL�T%��0�yi�*�����4��y<���C�d�t�_0�a����tp,�^�G]@��ֹ�nr�����@�j9)��Ȁ�����Z��}��ԛ*�.Q�w"� ��jyȰBlq$LahWV1lk���jE#�|IH"I!]�;�wm�%�u��ԡG99�(u�9ss���޼�Ɵ��p.��0�W�r�b��b��ܦ�� d��\-(��-�� Ca4��M̂�s$W��F�sVJ]ߧ�6�G6�Qfw\;��8��kP�:pۺD�qf��5b���FTn��*�dݫ ��Qz�/�|2��vvp�*u����K��/�7F$൙4#�<]����Sl�=��s�G��}A}���,Z��#������w;�潺��Z�{=�x��}�C���hgSC#m.T��x�؇�G_�"=v�L�9�x����z�>���w����Z��?vv&�-�'$E���LpS�+��������ZӦ�P��s�x๿���{#/8�;������j�D9T��Gj؎��|ԉ�+���ý.3`y���&ir���q�L弈�P��-l��R�2�ہ��(58*F[M�j�!�Κ���U�ݺ ��nc��e=��k���h4�0^���ܾ��8���b�~Bq��>ˏ���f�ʆG�I��\�`�s��C�n�R}3FnX��θ1ι��衁���R�%$ե��<������傝w#EG����O�E�{��Eڪ�Yq��r����9�8��2�ö[�0elQj�N,�X�7���I�6�vo�#6=����rs�������B%��;E�;7�$��|�07����}�SjY{ˈțGuӮ�awt����9���d�r�-cx͂D޻���c4��r=��7t�^�#�1����={�@��v��$p!S�*��4�H�f��5#��P���/l:��>;�7�H���5��Isi����<빛W>%Ú5��
�Z^ <���^��"�ind�=��!cCTҺ��q����	�wŒ*t��M���$���H{�Y�H�f�-��'u1+I<o��dqG�֜��q�VӖ�*��o�h��1N�Owo�t���)4 �bbd�Ɛ���,�s1�k̳27����g4�R���e"�ǟO?;��K=P�Orod�R���I�*=M}�s�V������JjB�ڍH�%.;l7��ķ����OgjǱ$�6�3Q�j՜D����h��0��\oZ�"�홷=���)@���,��.���}�LHm�wl��3��қ��<!M��� I5t�����h�I[RF�ݠ5A�P��2sﰹz��jvN��uv�� �P޳vK3��=�Җt;����1���~��J-���,�n+�L����ZrAX�������è�^��x�&Ms1�f���ǅ��Nҥ�Uϐ�[�I��qp�2��K5eu͙f2�5�ݟ7�p���wn�$�n�ɔ$��wu
)r�?>><x|��3�T�mΨK���XG�ci�7쇘�J�ŌK1�j�φK'	��VF7Lu��/zs�rH�#���-Q��I�3�,ݱ�����m�<����n�5�Ө�Ph��K$p�[Y�$Pg�T�E�)6!��P�A��h?�|I �3�st�u� ����xyf,�7��ƏV��\g����]���L��П{F�J�bCu�:�q��j�<JGm5�i~o�Aam�M�҉�~����'��vg�8�~	�=��3D�;���RW)�֎��OF�td̼5�J�=��Xֳ}�bEDiE����L�WD����x�}~>�y�����+�~zmc��#R0�AK[
��U�A4Ya����^��:k��3�Y�T�� �]Gˑ�B�y����=%pd�~�W3�pӓҗf��`y�r�U��黤�~CT�۝�j�O�99��zX���;�lU�ꮕ�����h{v�"O/k�;r��v=�u�9N���u�r��v�5��Y�l�m�1�{z^;6���x;���	14$;��s�%�����Yy�,ez�,ؖpC�]�NX ᛴ��6m@S������� �r���ɡP�!v�����X����kg�F�0x�3�M��{�����05K�%���S5U��G)��k-ѧ��s(�P�Dv��{U�OqyL����+ʥ�%ӗ�����WD2�d���a ��bP��|���ϙ�N&��E�`���u�gv����ܤE6��Y���Z!qh@�x_`[*��Ź�k��G7��&ȉ�O��+[�E ġК�y��x��"#/���8�"��E9�m��g�}��}����Ɠ۩A �F��Q���'���{��ΨL���^��Xǖ��B�H�*d��ʘK\�����RMsƚ�����U<��Xb��b��'�n�G��=��Hx2HN�Л��+�T�0�oj������iS��+4Fl��?Xed�)���yy�S�U�/H$|A$�|!���<|���|��y�=�?�O;:߉�X��[����-:�CC����J�Y��c�{��s�@gg��k�a�x�GbN�8�@܅�M�-7J/��j#�H����;��`��g���ta�h���66cԉ|!≊]�_���5�wxߑa
�d����K2%༗��C��E[��Lv��s�e�dT��!z!�+)� ��s�ó�A@S�)��<�瞾�X&��7�G�ۑ^)����o=��7ow��v�s���WwD���-�	��ױSܸs�!����t��t��KfxFC�E9|D��]T��Y.�wI�D^����u�j�8'�zF+k�:�KnZ� �ރ?~ǝ������6q���&�(x`���&?k��)��^<�g��u��c�d�S�����sn��*I��.]��@t�(��˛\Z�nG�K'k���1�^8ͫu���s��gϜm\W�F�|�;W:��v�MJ-�������Ɏ){]�3����6�F9�����jت����B-m����d��n�_4grX���v1����*�����;�Cs�OC���%�\&��퓶�6�f�Z��d�B.���&�����'Y)TuD���*ɬnL��usv�u�i�v��	�G8s�М�n�^���/n��\Bm��X��g��Q��i�X.K��n�M�ӎݙ�ɷj��������	�^K;�
:W��6뒺�ֺ�.^�\�����;���w��6����v��h����N7H4����}M�=} ="�3%�ɤ|���\0�iy�W�
E��w&��0� �E�+�l	���'��/9v��>*��.͖���f@Ɇ6U�/V��$�{{��G�Ӱ�z.,v��@����\b��\�3h�Qg5y1�EZ���P���8�n��҈n��ug��>��FzМ4��a�w	5u����K��F�SK )"�%&���cm^��:���J˭I�Rܸ�Q�jg�$��\�M�*��#o�d?3 ���0���C��� ��N�D+!^��rv�H�(��n�2s�p�U�خ2\�{ky^��Uʥ\���v�v{\r+�,x4nh7�w���٥��4Ez��w�w�Ɂ�\u�r7������о�
M���Α��h������W:*(��9>&�I����� \'��xr7�=4r�'�GePgfI���c,Q�Gu�2��My�<���rn	�+�&��]�w��C�_Μ�-��j�wQ�y�#�ˁN�$�		$�J=�k�YԔ�Vi�o���e��qh\c��[˅������0��c�&�Vș�(��*��㶧
x��7��g�h��.�G2[����v���MKrWKX^�m�^pe���*���3M��"�&����<� ��'����+y���g�cI��|�Osi�:Q\��8�S諢Q*�9%��7F*���+�ׯ?5vOw�w�[�o	fs��L�q�F|wL��t�qgT=�Y�Ca�#=����������j�뻿�A������{ݤz>	��@5g���	�ag�W��i�B�K  �
�"R����s���GA�*�(��#v}�'���/�=�aK�
RV������3m¾wX�;u�>�8#�I�EJ�Q���0D{Ԃ��@�O��1�0i¡�WOMx�m��zPψ1sػS����%ɷ\��psͣj�^
�9��q�a	�p;�mp�쒛5��}���?{럮|��
t82��ıp����w�����:tbM�B�;�HO֧��Q�D�n���8;�����=�7WZN�:���#5O��lM�8퀂��Ed��3�vxd<��w;�[����w��F��x:s�Fv��c��~����6E��Ă�>:cIfs��@��y;�6 �xZDx����r)D�����$��O�{RKG(B�rE*�X�dl�&�k9=x���{:<\־�p��Xc�<礫d�֘�`1�����ʪ.^��r�;������fH>'��Cji=%Pf��$o) l4��I+Q���SqlP:���A���"� Ί#N5+i�+4�vxJͼy}����y<�"��6�<؝�Qr(x�;Q0Q^�!GY53�����Cq�V��=�W��o��>����V�(�1�@O.�Er������G�ޛ��gN�2,ECZƣ*��P�k�#��|��J��nb�h��xz�.Z�<�3�]��i�M6���fx�g1~ �(�� ��y�1���a-d^�U	�Z��M����g�C���a���`W�?f���հu���K�Wr�ǲ���O#�COax7$�9��ۦ��"��8�i��vhܫy���j�Q5�?{�87�o���4���e��D��:e����7�rMo�̭��=��<�yA���G9�*�4W��gH���z���+�x	C�}N��=��X*
䎶T�J�n:@,�JC�X�w���	��W�;㝚�(F���$^�P#K��/�Pg�S�Ȃ:RzRl{�:
mO>�Ǫރ�)�׽��𾨎r�6M	��h���lG��44ݭ���L�[�ʣ�-����tu��V>�< '�[pr7�B
M>g7Y�5��K3�7��t�O8sRz����/��x�qh�\ޠ�>��nORf�A�I����I!�S�3���ڏ����a��5gۑ1q��Ggp3MSR�Z
�S���;�f�3$��.��'2���C�ڔL��� {OA�{I0󕘚���W��^�S���sG���{�:ג���po��^�{����FJ���z9�{C�9�V����g���!�xJ��{X����M�N�M�A<*���c�	�Y�˛I�I�̧��ygA���[Bg(����2Z�3��Tk7u�Ypʭk^9�4Zؤ�C�z©+�%�FX���m���#���a���m���_o���d��s!�|� yB�S�3Ҧ5罸�������|Ҿ4��2 7R�Y<��M�'��_IJ����@�>�S���"E�j�d�^�ǡ>׷*����yv����#���15�w|�#���������dYd�A�#K[�F��,ʄ�F�-vQ��&���Y:���!�2�ٕ��n�;J��e���b4�I6ӉO]/��Ȁ�{�a���P�ē�}�ڟ%ӻ��������+��q��w���������V� r� �#j���m���x������vH�ߣ����n&;F�6t��âV(c~��R[�ׂݻy{�o�aZꌙ����N�\��j���|$�3�;��L����^k�����{�[H�q���ƉSN¢k�3O7ﰧҪ*Ic49�:f��6��Gr�W�E��Z({T��P<�ݣ�Y�u,����ɬ�	���~m�FM���,d��.���6��&�a_-��,C��#�A��L�����e��|����^�`Q��ӌ��\��ojd�gC�n���p%�g
k{mʵ��������m�jUykj�Ƭm�ʈ���kg3�bw"Y��a�0H����n� _���v��N��#H�R����������C�-=��ݔ+�YY�9�+,��z�C�X���l�"�L��]������J.��{=4��h*Z����ҹ��F�P۹{��(2�2v���4V:d��>�x��,�P���z��0:Г~��XW]l�C�l*����K1k=�O���x߹p´A�J���N
֘��4�)t4�1���ڋEr���b@j�ʒX��w�#Cf�8�/�k��������z7m\���ʇ0k�����)�$Ѿ5T�u "�H��4�.�r.p������H�r�FH�"��UWk׸-���bu�z�<��=�/�5kec�1�)s��FǺ���)ݢ��ƸCK�Ѡ�)��݅3�y�Uʒ!��Y����.M������\0�[
E�q�$��.�2�+p�t�#��Wa��>�0�-�9a��@��y�Pr,ǁ��/��e� 2U�ǩ�#���P=���]i�)�m����w�4_7L/s�Ip�/[D4^���ՠ�h�)f^�tS�X�y�em�n{e�9�f�\X{yֶ����dn2.�I����c�ͮ��û72p�k�X���z\;cWf㎎������}��W�
ah��u��b��k^2�{��2/���gڰT!�k���؋Gbc`嶭�)	,f�<DB���:ٸ3@�[�5=�q�a{�/�j�8DEkNDr�S����:aЯT�4���c�}y�s��t�Xhz��\1��\�b"���7IĒ||O�!J����n	��^���$&�`X �+<�<1n�3��3�.W~L�q?��$��A���;Ik��t�^��O�gz���4z�.�uT)w��	�4���^�י��7:��b�qOK%��]S��ǉE�>p	 �m�0�I��k����!�8�c�	#]5�����E� (ʨ�H��RW5�R�0�\:ib�#o 򣕺�ä�L�jM{�H�M;�h�����a�	�.��N�����Kճ�	�c{W���"b�j�5�$�Ĺ�j�T�:ױ�e��4���{�qJ�DF�6Z��ڪ�T&��5���B�[W���D��K!�m�+�b��#^<��?j���4X-�[
F!� .���g�q:�;9=`�=Č#I�$�I! �QA��
A�|�4�}~��8�!��5�9i���xfL"%D� d X�BةDIm4���md��J��[Y��[s]���լ��e+m�j�j�e�V+[FڨŪ�V�r�[�V�[Qhը�M�F�`�F��"�j -X����Ѣ1`���.`����ch��*+T��+sTmb�"�X5��sƪ��F�b�Qw��<Uo+[P$@�D�Y9b �5kՒ����Ѵh�Ʈ��6�b��F5E��Z1��Q�X�TUZ���mm�V޽zx���m��Z�V�QUh�8�4(b(� �ȥ��	�ڶ�kV+kĶ�M�b+*HU�*��#b �l��P@cRA��1LDA��2*��뒔��8�4�;�Zf��&ϢG� �+" ���E�}�?�����>�Q��ާ���~��������w�C��y�;����_����O�vd,�=���g�M��7l?����=����?�c���~P�}��	�x���A E;���F�����X���|������a�B��_��Eo����O����  �A<bz�yc���O�#��:0Z����~=ပIY�爊?�ņZ}$l�K�>�|���=�h*(r@,��kL�M--��Ե���Y[J�Si�J�jj�R���em-�֚�ZZ���Mi�M�֥l��VZҬ�Kf�-M�-���miVmi�������Q""�H �X(�B*�D��T"HCY��+YKVSV�mR�e6�J�ZR�6�l���JZSiM�R��6�VR��R���)���J̵)m��JU)��ڔڔ�)�JkR�lͪR֔ڥ5e*�[JU)�)VR�ʹ����Sj�ڲ�Ԧ�)��5R��S[L�R���k)��[%����[e*�mJU2��e6�-)�����R�)m)�L��ZҖ��R�T��)�Z�V�6��Jm)��32��))���JR�٥2�JR�K)e-)iKJm����3m)[4֥6Ԧ�)��5l����T���մ�mJV�-R�Jm�Ք�)R�JZf�6f��jR��L�R�4���)e4Ҕ�6SiKJj�ڔ����ڔڥ5���3[)m�5Jm���kJV��R��M���@! �SL�1�\A.֛7|�9����v���ߨ ST�QF�B��I�{�a�?0��Ԍ{uǭ��=��>��9�Q�`c�|F���8�ϙ@��47�<~?����=��B�_�~��?9��,���C�?G����j`>p�ǰ�����~G�x�A� �o� ,I��}@vO�>C��u��;�&F!�Y�|� �ϕ S���Ҍ_���O�����A��(�C����:��G�@�"�����o�DN��
~m }����z��@���c|0=�%��A����a R\����P��$ O`��x>���.����}��~��1�C�p/��C�a��A�_k���	�(��3�:X���G�@?�=��� �yQGّ���=�O���'�#��#Ճ�����S,��{`{���>��>�X^��w���S��4�)����qEQ���@�>�#c�@Ѻ<@�@9"��&m�<���}yP������)��!����FOO��f� E=G��R(��>֗?���i������?���A$	�������(�g�����?�����]��BC�nΈ