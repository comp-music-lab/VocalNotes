BZh91AY&SY!ےz �p_�py����������`�?�         9�U@(H
UI���      
� ��� ����}�(�,�t��.v�)�I��r�KA�>��J�U�qH�����s�R"$L��	$�[�W�M��t��7Q%gY�"�y��T��w7�QE��(�Gs�E�ҷQG�����iE(��B���
�<�(��vtQB����1�G�w(��.��EQ꨻�P)�\'uoQE �gE �ugE��(�YIR�g(���        �� T����F�4d� �d�h��D�J�2 �M0&�LD�*�Ji�=C@�A�C@2  ��A2�J�0�2 �&��@bO�JI��F& �� �L	� D��h�4&�S�Sҏ��4���6��M�j�ǁ�ǗO>���4k�*��P�@$� E�������P��X!���@#Q>V�%T��\@f � >�0PD)L]#��l���om�DA ��B�q�3�)�$�s�I!��+p:7���2��HT�X���/�sƯ�sI�M+ӣaҐ���j��Z��� ��DƦ�О��/z�>cl��e��ټ�=��F��V�'����{u3�f0K�;b�u��̳f�bѢћ��x3V\���:C�ܤ�2�1��:�'�B��� oN���9$zm|H�}�B�9'%nuUwtY�uj���'ݲ�٩����d�3h=Ǟܣ�Q�VvC�	:�t��ӹvq�\�[�ܸD���wu<��7@������F�W12�́pJ�g��(A�@����9r˴)I�Gqk��;9��e1��Qt�/\Dn��
��o_0wSg:�u��l����G�/i�繥�����5Bcm^ЙUg5��O����1���O��:��G�%rkf�FGi܊�:A��żL��u�+c��<ԧ%�i�(� N�SM��MZKZ ��5��{9����_�6��F$�f���K��P9FD��8��9�:�6>�ۣ�y,3��s�gD1ȭRj��CX��7�r��&��lXn9�2�cw���n���8j�)�NO���o���v��F0�Is�����G,�&���;�.����|�t��Qtm�Q}�сB]�pzE�{��n��\0�P�"�ӳ�s�w>�t��G��8�F׻��6�Mk,��d�ˎ�����'&=P6s�`zw��5Q�F]�S��3�\z-�X>(m �h`�CD���6,�>E��Zx���Hѫi�9M��Ր9�;8�v!���7x�)d�wp����6�l�=nrÁ�'-i��¤�%��נ�᩠�Z�LoE46��QknwN��x־§s��oG��)橌����gP�,k���L��^B(\�))��h}�Sr=ueY�n>��z���+�Gv�q�F����C�C�r6�]N�Y����Շ��]1`���0w��z���{��ݲv�V�`�6�Ά;7w�b�'s�X�����9h���K�sQ�_�	,�]u�j�)�w����{^9�C��9�O�фok{�"1�H7�t����+n��.�h@8[�n�l�+Uٛ�O7�xش�Q�񫐯���gz��u�)���6'ؕ�zAQhoK�`I�ǝ�Z�*${�'��X�{�����gL.-[iX�c�����'p�Ix{����!)*�yk=F'ٷVB`e	 4�o7O9&�bEV-�\ �
պ5�Yݪ��h��v��e�[����U8v⼖. ��L�(�~��N=��6dJ��}�v�3{-
c�N� |�[���Āĳy�o��\��۳����.�.�;	:\�����B��e��sz�Wv��-�'CwS�P��I=g�Y@��Ϥ�.7nhM���HK������ΎSqwQ�>��X���ůE��`ޚq�L9��H��p��-�11P(��.�W3xظG �#�H� S6�$����V���/96�ҁ;F ��N9��M�w�0���2ds�����^�5���5�u��n��U׽�^�tZ�e�h��ٱԐ��t����z���\x6,u9�����
��4�v���Y�m�p�C�܇]�e�1�#9=<a�8��N�ib�D�����E�w)�7n��UB��U��nh�B�2��������͏@ι�pȮ�2��|�t�{�m³~�`a���qh����ݚ�ם�1�����T���v�3:ˤ��p��X��Tn^96�9�d��9�F�E�s�����:0 �X7s��{���r��K`Cah�2[��iH���:-���+	y�T-=ܣ�h�z*'�ɇ������ %��ܸ;0a�t�X��klOo�?HUu��ʧ�3��ɢ�C���x�:6فQ�����:C3=�^eG=HZ�{���+����sn��jqT:�:N��'.4��nY�6��V͟Z�tץ��Uia*3:\�S:Y���wK�㮩�嬻U� r�jV8�b9���
�.DSn����F�:��)�Psm��{x���$�@��]�=^	p�q<���F�\l�f�!�Ќ�M��7�շ�庴+���k-{6�ۂ�:��gL�`m6 �Ghcd׎�^7]t�6B|v�4�4X���/�,ҷ��&��=6:�g�]aWۄ��kh�����Ʀ��f���q��t�:cq%�]�:RiGf�fY9��ts�筅o:gyl��ut�W.\��e���k� 9G��N�^u��z��с�����mfNc�c�a�]�5e�m�8��x�.�*���`��q��X�O0vc6�m�5�p��6�]�;E��ݐm�v��Gi�i�U�`:�n���xѶ���f�� d{m:�ԙ�quQ&t���cؗ�/f^��ض�d垃���I��u�6��7�fӮ��ͱ������������1��8�π�I	�����n�{��<�H5��d�[&ۈx��l
<\������ݗ�ZY����۱����l�Q�a�t����A��VZ[�z1�qљYL=�l�� bg��vw/ssx{�H�����랻K�m�v�a�u&<��\��V�A�.u�u�&�룍9:a۞kbVW"���x��P��11��`GC��U�hMn�oV�[��Ls�|����=�.qlx݆�s��.ʞj[Q��@'Y�v��N#Ӟ�s���3d������p��Vmy�Tt���h���n�M�%��%k\�^Gq6Y���RQv��Q�oGn��\<��1���z�y�]�<�vB������������R���Y-�Ӎ��8v��ժK�Y�J��QWq�95	p@�efq��Nk��-7��U�:��7��s�;Pgu�u��Z�d�v��ovy�v�$����V0�7���ۂ#ۖ��E��ikl�8�ƴN�gL�"b���ؘ��C��n0`�S��pZ���I�@�MZZ���q��GE�)˔�Z�Uv=�q!�bۂ�U���U�t��&���-�*S18�P!]ZR�&K�si�#��.�ݷV1<<��=kq�عf�Gaew�����w7)�Ӈ��q�5�5\�S�.ョF�x�e9tK�n�a�G1W:���u!�(��Fx��S�Ŧ�P\m��� [�u&��뜵�M��R�����m��G`{\�"{y���EUu=
x����]#.+=n1����]y8b�{;�&`B�Q�rF� �|�v�!ZUwXlN�����ո�b@�4�T�@/�<�N�1|�z��}9�6��~�[np�}/l��P��g�̠�Bz��)QaSvr�O6yRg�L����Gv��]��w���9�'h��;ѓ�_xyl�I�ۛ�v��ot�)}�.�Z7�r�#g"y�p�_Nz4�Y�=ڗ&���Y{�yY�p�^�tX�a#�u0.
�tS��ww!�F��������WW���M�5�p�E�%6�ܫ泊��Vm�"殮�g!��3�{��I��r0܋ƽ�`�YJ��:�O|� �]dvh��l`]�`x���f�1�K����z��.���6=�53���0z��%l�������ֹc�v1���Cݔ�tS�[M=��A;�T�|������xWx��p���iЏ��8���O�l{��{�����i͊Ӫa=Ȗ��-�j�����w&����8�;�@A�|�0�jc
{�����qS�G�x�ޚg#���燋�5�c������xh�O�x�n���[{:r�x_\�eY��f���2��lrD��o��c��vr]،g��7������4�{�QFv烚bX���#/��}���#��VߴZ2=�I�⑝P�nw5��Ż2J�m��Y�W����;�s�U���!��2Ozo����O{2T�eO�ģ{����}nw�;���a�s���=�"�v痯�_��y��ý�}�A��n�Ό���kə4�Rr��r�<���Bִ}�<�����dK��Ə@z�:�W���'[�酏g��l`j֐��C�aM A�%+��U��5{�Q��'�LXw�����{�=��.�<���Bf�3���qV��T����y?b|�8�6{w+w���:�����<_���k:m76�{OVt�F1�}/9s��{7���~<���{7�}<zD|�vm���7O:ǜ��2M�����Ι����H�x�`�FrXc����a0=���HV?}�O{l�	�A����"��N�:މ���p�Y�m����"�l�t:c�l�7|�	wo���N��ǯϼppj|�Ǿ�g?�$�N���b���gg��°^��> �
8�ԏ�H�3]]����!I����CG�k��j��E��vi�A����w�&���|�����\K M�j�o���&��G�T%�[C��8�\�z�/��c�U�����t��wP���zR-�p�=�߽��N�v���9�D���m&%��WP�;pm����Y�ń�o;^��g�~���g��`+}:B���a��s��gx������={=i�N��_���`�obTX**i�c��P˅�"��5�N��v�<��MK	�<0yv��n��6a������0s�w���
�!�7ǩU�gu�E�X�v� ?d��K�Wgm��m+�v�$ml���/Ҡ�*�����=7�o����O��{��Mx�W���,Â�8^�@��6�&�w6��=�벾�b�g�`�|�SO9/U`����]^I�٠���`�[�9�f�p�8��/�������s�3Μl�z=�q��	2����L�v��=���5�rm��ŝ���v{X��i������7�����vy�n-�B�n��C�t�e8�2O����U�x7��;���N?zdٞ�̍'9w�<��|��c�s\sQC�͘��|�zz&q�W�_}}��|���ǐ|ТQ��=�$1������}���a�V�g�~����p�2OS�7��7�w޷H�����gO�x�S�k�ΐZ�vS��~{}�MQvA�J����ykU�^]�(ۦJN{n�:<�6��8�E�/ {����}�ŝ��������|o8��ی�����lnU'8)�)���MC�<��oL��&%���kpBx+9_G�7-.��E���g���s?;��A ����y̾��A�%u�t�{�|��y��/>I��㒙t5��6��ռ��i�1��c��7c��R�ˡ,q�x������י����l��Kr,��;,c��T��,��ьT�c��&�,���S;u�b���뒎5ܐ����Rj�<�뱸�'z��#Rp��9�{K������GO���.gB�VD�uZk�ӭ۱<����;G<(7��õ#�F�u���^mE�FN��9�V�C���We�^���J ��(��M
��M�cvJ�2����n�{'Bx8�S�ݚ��g�.-'g;�~.���m�ߠ3��pm�-���2.��F� ��Uf�-ʤ�
�yN������l|CW�Q�p��?���^ 'vy�ÁG�xh�����P��� D�@�U�5Bi{af(�P�h'TsY�I	y,�������I[!��\6�al3,�-���w̒<�YFJ�x*�+%� p~#����P��5WT��ﯾ>Z�|�?�E�1���e7���I�6�6����G&@%�����M�5��j7E��������DlCr �87?ۊ�̟~c|��6�k�lÏVv�gw�g�7vC5:�5�bo���x��as��Ik��u28��:>L���(̿
֤�dSe���h�8v"b�M�Iܵ��g`�l���zsD)0/uk�	�}Sn���	Ƨ��NN����W �v���,�u��,N�����N)p-��l(F�6D�Hy.�s
��s]�5��P_:�A ��Tw�����V����^�+��ZKr�ك��RƮamr��{������3;��ӳn�T��9���^�*Z�Z�諼E�k�a;
r��ځ.���|T��7z}E�ʢ��!���;d:��g��Ů|ۙP=�I(Y� ͥ��Q�,��hkl�f�%����c�la�[��M�ϯz��7�U�m�%��*�p�c͎n7m���L��:t��8�rwg\q�D2���;q�sby;<�|_f��U��3�d�ݦ3|*�z��v괰�j�$i��I�{0�^8��@3�Txw:�몓v�������O�ţ�]�9�L+��X��R�v�8w�^�m��AU�T��cכf�NŻZp�O���]k�3�u<��RZ���&D�r��堺�m!i�w�{��0�c�K�i�	�#K���s�sL�m�1�6̛� �J�4���{Ԭ�/�CF�5�]#�W����AZ�*$�4]�Ldi�4ٚ[�ݚ	C�5�k�"f��Ka�IH �p���`ȘO3���oCT8�,�!;��x���5�R}�jvQ�Y��"��V(�Hb3, �v 햁^,F.<�ٮ���Nh^Ś�<O��ap�vmؼ �"I�ֵC�^I����9_/.l�O�V�?g���D�n[Q@��Og��M{�ܞI��s"���X�[_H|ם�	�z��5�f)��kYm��we]�D�[- Ye�ey��ﰈ�������,��4��4�@-M�����ҵ�%�>��Ao�L8!�����p@TC_|e�1޺i�;����v6�i�dҖE��[�<�9��"�63I���k�I�*���e��_=��j�>֧H�:�*�`�E�NE#Im8k���UlA�-C���P���Uj���*�Eخ��w�m=��jÝخٞD/��٤�=������ǘ��M�:�ϷfpJ����	v�<;��RgR̞F�n>T�RX�B>�݌�-'r��L�������%�����o��bb�Mt,�3%��||u�n]�}�2�[��H��֯)�mb6�);e��Fo�����р۾�Bpӈ���5��g�q ��6��c�u
B@��j��/��wGN��ppHi��-il�\;�p p��γGP��z�#��u�wu�yA�^S���ݷ�`[ UK����, Sʷ��E86�q,(�>ڗ��f�tVA�x<k,��^xr�������]M�D'�ř-�#|#M�6Y��7��oň4�c^:g1������,�f'��cĞA`�c��c>�s��*ep�#��X'e�Gu���.b*H ��lwh��x(�>DE/ �v�PF��.�i��+ڰ���
�z��4"�h��R���Z���a��| 1�>�䇁𫙻\�����\dS��v�׶���>��i�� k�D֤M�v�t���1�٘���gp� ���IY�f+��0��mm�*�� �k�M��e$5֓0"7��J�^5ΨpF���*�]A�%@6�DЊ���$3Ґ���^��	x1�6�gT���CAC8��n�ݦ׾��iJI���G��" c�}���y������e�ﻧ���SFn��|��:�Jb��B���j�q6�Q�4��aV��b��i�	v��/�7D�����g5�[��u�1���D��rqf�/y�C|B�̩*�6 ���9JHo���Z�b��K@/�n�C8��h���n�T]Ѩ$���`�Pݺ��"T]���ڭ�(� ��$� mIP0]#h%���ҭy�$7n�-R(e�o��TÖ��I�r�(��Q��l�XR�nvߙ�~���ى�f/��kC0�Y�V*�mSי��������#i��q����y�i�>��N$񄱊�=�3i�� �"`�H@>ʊ9��ݙL��4���<`�{IԢ���SQ�CX�I<��w����ϰ��0��t]3�J������G�xE��1�����S��`H�h/%D�sf�2iy�~��� Ա#Vaq�� .g���Mc�#��Y���q<c��7�g���êX�,��Q�,a�.]�OjY�g�b�l�*� �&��{fp����Z~	�I��1�>qm����F
=���5A�tyK]�U���xѿ����<�h�˙O!$�K���<�ּ�a-8�#��6�w}$��� ��*��KKey}�A8$�H�o%�2yg��yH�F��������+�%	W�|=�Aot�;���ǘ��XOI+{��-�~ņ�1�`�#E�μ��S��M߄1�U+M���U�����ү����T�GDo6�8�9�Xn:�5��v<��(�i��b-����O���#(��U,a*��Y3�%�:��O@�$j�=����񏽑�KX�#�y�"�z��K	G�b�X�ߤ~Xi$��h8��I��~c��=ag��HUl� RYj��KJ3$��))H��ƐO�{�O�ue4�p�˦0���&�=v�;6N0>  vc�2�� 
���A䌥�D������ָ�cǡC���X6��;VzXx�0�2����X�4��- 6[[vQ�[u��0�s�eO$a#�<{���O��m���l����+�P�c)&��,#�����txF�H�ī�ZZ�����^H���S/x�{� �G����-E�� S)H�Q�� z�.�gs2x������Ny&@�W�z&��
��)U5�,a�\���.�� <�(��+N�d� =�{yXx��#�RA_���O��f6�=�f�{�k#�AE��9�v� ������fm�  � D8���O���y����ȽU�Ye���˻~�~aD���#�����[��=�ILa�oc���KX 9��i]eW��i�4Ǡx*!�y��8� ��Q�a����j�!5*��W��2�����*蹅�I}���C0kɣG�������{W�y�[3��V�g�-�pw /=�P��3���g6�V_WE�#Ӡ�r�r�][l���E�1_l����݂��= Wݝy%�y��|w��=E'1X1��U�"���n�ւ�c^�7"�w�����S�˶,E9%1L�Y�Nm�u=q�rO{g�@����;�Ww��T�d*�VGi��`�W�i��Cd�qۻt�f�p�l�Z��=ׇJ]E�c�ۯ�f�.83�N����N��ִ���ti*��X��6Գ�NY=��Ų"�=O��87�����v-��g�i.!_˙��)}Oϟ8燔����Ƙ�\r�ڑtAcwn6�ǝkJmw�6��� ]�cs[ۈ���T\��GvNݬ)%���-��2#x``�ep;��g������Ӧ6��6'Uۢ佶��Lg���wl޽=��k��Q�ي�V�loX��N�M�Ŗ@^�������b޶'t�u�6<���=Z�諾޷��f���HD�Y�MBx�s��T�q&������0�<�h���-6J ��Ut{,�&7��tEdO�.F/�D}�Orog��O{���x�ۛAR���z�_<�Y��31q��p��Eۓ(Y��%c��r���ۮ:)��ur�˶�*�v���������PF*(ʜ���29^j΅\w�,\����;L�Y��#�+P����;�ƕ���#�ǆ<��`�#�@ʭ��E��JV�GR4��27�ܔ�c*�ׂF��ۙkޟ��~���%�j��&�W˧j���L��]Q�c���6����y�;����H����t����{&�r�6�Y�A�c�?�e#��$��D·mQ�X1���#�N$��?{Aǜ���nH�F��κy'�QIJM7̖T7D�#�[\��Ö�S3�.�U$|r:�ml��ƹ��M,ϥ�ʃ��S��yKK�]^ET���iKUvK.��<|�6��~�=9�)�>�G�%&}�yY�xN(xG�x|�;H�l4�$�.J��㬵�DV�O0f���"N
y�h-�mHճ��匥2v�5[�E*���ӊ�{K^����;�~k����-�~E���lv�k��\��P�e$r�ޡ��f;����4�7��u�Ҳ���[So���y7�h��l��,��t�b�X�n4uݔ_=������ڲn�53}_�κ�u�����VT;jc�X�3��ʹ�����QY)�dy���}=�9����ߦ�)�6��h8���aq���s���Ԟ��F�/W}��ׁ�����3�c>�zR��lTC9"��IԌ����jH�o63̞ɚ�&�c>�e�K�|��K燽ؓ�a_����6�5'J�뱴��4́��@�#+�{3��}��%�(lp���7�TV��DQ�E(�;~���2�f<�Ql/����ԍ( ��V3����&w�Lb��K�&�6&���^��X��Ǩ���t�)]�ygw���20�ԠS1�<��̞K���6��{z��6�c��G5�԰��C@���)��y�C9�q#�~�*z7���H����${�[�����/�ɾ�M�jd�߫�>��-��f�&>��[�c�>�،�-�~D��X���lnK*�۽��#��RP]ʞ�2�qC`Z��>o63��{Ô���x�M+uO��~�MoЇr����ϼ������r}�����jV�Ŷ�Y+G�/b{���q�̛vw\��BV�͙�0FA�]ZK���H>��K]�w���0t���K#�j�_�|-���o��\��<�[�Z��E�����&��N3���h���[����8����J� w]p�\*�\D&E]1\-�Xo��4��,�>I�z)�<��e��R���Y$:)x{�L)� �a�f~:hҨ�E4���,����Ⱪ�U�>���숥�:�:5l��wǧ��O:/���<�޻og
�1�L�D>#Q��I2���û�N�&���+��(�
��y�Ͻ�
�7�YN����;.Z�˭�|���'u[�o�z�sp����g���x�ӞR�*l��%��?$v�G^'~M�_�J���T�9o���r���Y�qW��_Z�sݣ���:�Y�vw�|=N�y!o	�jj��:��ǚ����7ӧ��3�{N6N��iA��1r�[�XKPf�)}d��z|���1��0P�س	 �Z�%��Z�t�	�z���=U����EF,x�s{M�-�:�='E�j��
Q�*�3����a�1#��+�	:�m]3��&��"��5b��22�x=�����Mn̘�d.1PL��c\5Dv������U��֦x��oB��ƛ-����;�#�-MH㣅p��yֻ߱����L�x�XB2Xk��27S�k�t2�Zެ��X�;+��Ю��.�v{��zn}�kθu,�a�������V����Br��[n�2|̟y���y^�Z�L���^�or����5xf'��L��hW�2q�S4*��×){���lѭt���ｄ�VR�R��� LR��[[��9�r�v���5��TN�3��ց,�4�b�!e�7k�GC4/�9'8r����[n`���]���g�pW�r�g��͝�6��\���B=���PL,. ig�]���A׉����zQ�c��TF�C1A�犅�����e���arǳ�b��XY��ٜ�wۦ����J�ʪ�<v!~:�z�m��K��Ǧ�t�n}3��Dy��λ�qI*r�h�ׇ Yl��~.�Ę��nzٕ�;��-q�\�|J��WYCa���w�ymSg����yԐ�"O\=���T�m�񚓻ǽ�T�Y���MPRWZ��b����vY��ۗ>n&.:|5�[t�sE�5���dq:�Mb�I�%u<�5Ee�r�"�L� ݰLŨ�4
��BUk�x�Uu� P0-�X'h)!��Oa4��#�<�fZ8���Vu�
�x���%���Ǩ�ՀM���/�_C�v���T[V�d)�y�b�ٖe
4�*��.f3+)#V"���-�ѤI��s� ��v�	�l^���)����M���*�ō\�)û;vx�1k������z)����jwh��^��mS�b�<_�b��_���ދ�Ky������I"j�YJ�&�֚��So^�O�6�n�ܼ��-U�ݰq������a�Fva1q��-�b�ץq�&�n�+�u�sqy����R��+j�idT�5浓��&��Nz\�|����-�Es�	�V-�P鯩�ip�}ݪJ)º��|7V����g	h���Q�]%[<n����4\8pj:`��t�q��^�׼V{��/k�s�gW���pouc;��O*���xմ��W���q���![��u���Te�˗I���wy�<ˍ����0E��(�%�#V��4w��>?^3R^���;�@
z
A6b@&4w�����r�������hZD��k�Z^�3���d�������uŜ��ID{�݅�����ѧ�w]��oy�%-zO��a��ӹ�k:3��l:.]��&R�6����Q��hI��D{P�a��3
�p��˽���1�%1f��o~<����5}�<�����uٛ�_K(Pw]�#���}Ϻ��|�Ǻ�ہ�غ�E��Xgr���������|��t~w�v%�5���Ms/\5�{���99 �%��U��%��l�y�-�X��g�p=�>;<�.������<�sWOkv0�� ��ϙ[�9R��ng�m�.����.u�m�͋<�A��tDv.��F�&������s�u�0tg�ꣂ.�j�1���&%�R��qt�6���^õ�:G��[��q�a5���x�7��h2�J�k7dMy����<�1v7��t��L71�v�aZ�"#ܔ�U��ۯl��$��-�eA�F]�^l���eo�ܬ+Y� 5Ib)C/��L���x|y�M�N�N�}�;f��Kؐ�2�$����_L���1f�X��5�àp�`��d�F����2)����6-� 9,oI�b�T�����2�i`(��,˞i���3f�"��Hc�N�$| ���&hSf�Z�L=&��	����� ֶ.-]4�r)�/��wX�U��7����G\�n惃qǫn�WZ���2���n6-�9��34W��&�ORI	woi�tͩ+��Um2��tޅ��o�93� $x���j_5g3�ҍTG7�&���g��Ph�~�r��Q��R�J�"ˁ���]w��8�Tu�����f�K��:X���TTP�.����Q�� >�-)�w���M���P�[�8��,
�C���u[S�G�-%�޳fRW��D#�D!Z��6�;�Q�
��,�>�u
���e)g��u���v��vzp�����T{��Qzr�M[�(���`��XOpZJ��O7m�)Gkn�gSFN��۩W(�V �a�?�?��!���6j�g�:X�SW)�Rc��R�5�R�2����mnxKGhl��=.�g�nR�(D*�*�+5�Z���U�����e��z���Ƈ�Zi�2��/Ԝ�p��gs��L4���v��N5���
�f�oB0��7�뫚6��k	mv�����tše*P�E���p����zS�D�a�����/W,Z|��{�,�ic�j4UDK-��kM{�BSG���Z��	��.w�I`�W-���e&c�Ĩ�)�hP��p7 �,5�`Bq��c��b���;�)͊��x��.�-"9��6���<uχ�!�y4b����XK��n�^�!K�Y�Ut�],C�m\}��l%�b����NZ�2.��:�Y�h��
h�b�O�-�7P��ˢ8���;yX�b�R��g˜!����6a�����PW(�a��o�3��b�k����r��6��7�(4�d-�[�r.�����v�>|X{}jS��'�s�Q���ޢa���ܷR��g��.ݐ`�*0��T�x�a˨������7��~<!���i37;�̘V�IYk����Zg0m��z���ˋj�R�3���B��T�b�s]!�@e�������iR����	����|&#ō��*��W�·f'��#1��̕CM*r낅`�4��ͱ{^ۍ�͵u"�Oh�7gHkw��z��r�"��,V;e���,�^c�p�#�yh���B�B����K 铽�m���(��k_�Yx� �ܪМ{����bL S9e��}~�[�6��'V֮�	�24*nWV�C��|hbh]
�U)�wuC� KR�<��Ńŏ�7��f/��nm�1��3�Ik����q9+�&����l3�R	�,h���Ja�q^�'a\����Q�=XL[�b�Wa��P��vQhU>��j�����ӘU��ا�ܑ�wܸG��r�tOW�+>y�ǻ���N�����v���~����N�3Wxנ(�y$�j^�M�s���p��-\U;�����fz��ii�q�y���˒B�n��}�	��/�:�I>�Y	��ہs��fm��j�k�4��C��B�Z�`���Jݽ6у����g.W�y7�1��������ظ��~���,�Q��C1e8r0��&*OK�{�B�ö��{|gF���G�I�,&(99�Y~X���J�u��2����������a4e}t.��{b�=����Tq�|W��
����F�D|��#ֽ��-�;R�Z���kv��8���E@ �A�����Xp���O������n/1Ռ���	)!m(Ю,�r�d�ly5'�]��;<����8�w��=�\��4�[w�5n����{f��,�[fp�l�(Z�=0�5�����NRv�;�m�)G+�^�Y�j�;�V3�ߓ�"n{��8��2���c�Qn�B%i�56��\�eƈN3Xf�^<�9@������o4���J,�� �5]� طbSl��6P8����8�+��9��f���XF�QHH�=�mq[Vz��s׌�.�x�U���qh�>���;��
z@�b^LGt�d��{�<3>�t�x�֋�ui���+�Y%���e���j�CJ:�j�L_|�%i���S���fݩ��3�;<� v$�r�����F�k���&��&�7T�<��Z҂�M<�v�OT���nYc�+r�;���y��:��ݿ4�V��B��:���j�~�S�b=8��<�<�Ǔ��z�;+ۓ��8
ƪ_������+]�>�yo�J��tx'r��0pİ$�S����������~���'�u��-JL㌀wU�I��<��yp�,��W*:B�4��J��r�ˉ̹B���rz6��J�ɵf!>>��ka���(��7,�r����-�~~�y�0�v�G����hT[i�g��h������V��^�Nm�i��F�5I�� i/�v����9��7nrm���:�0'^��M�j�j�;nv&;;��zO7ET�G��K��c(��i��9fg.�G���ѮϹ~�����d�cPY5�-���֛��4�#lL�'9�mJ���;\	J'm�����O����l��I�޽,�J��2mMb؅,xfdx�'Y�����):M��w��氻�0�;��emJ�p�çm�9`]6QR�(�o�R�g& �y�P�2擾��ݹ�E�Nޱ3#�mR�cwÆ�lyN?�}��ho�\5�;�ъ�����ddN�מ�Ė�/x��6d��c��gܚ�Ԇ�x�s���TZ����z��\lY�m�l#[f�`����K���uɅ��K�B8F�����w3�`*ݩkw��8���R�c�'�y$�1�[���Z���}�n�&���SmM���A���5x��E�ա��\����e�f���.-G&b��mڋ{u��&�:�O����Xwy?TG�nn|�E|�2��Jeþ�8fyv��3�='�GPҏ��xz�n->��)��R�9tR�ІD|�Q�ȋ�x�cO��M�{.�5ؚB&�K���M!�dE�M��Hq��u=�w����]��8Cf�;���wp��C�ۭ��t]^i����k����r�MuN<[���ǌhX{�����N�p=W��q����]�Ƈ�2d��Fs�$ �R����lэ�3Ŗtln:�����lL+��If$�cf���-˦�f�-�t�7o^�dAa�����ڇ�4Aȝ�T�҆�6�㛍�]��Q�V�^mci��@I�����Ӎ�N�.Yxz�v#3.�ͦ��r�Li�^b$�����Z����G�a`�l�u�ک�m���c���l�9|���꒑F��x���(��Hё
�05���qEE^�ɏ�s2i���t�"r{[�3�0��h�Q�f))�� �����nh���xn�-��2�/��&5/=3G؇�%��2FtQ��)�X�Ցjȏ�i˧05M�<�I���hy����XO1���ѐ|[�}�hW� +�X��Sͤ�3��g�D���ᣤGێ�^Ą��:YN�u=������w��-����NZ�e�@��Vs�T3���qmYj}��f�<��v���Y��k�4�km�9��}���3Fq�sp�n֪*()�DbE��F�
����౞:;l�?Co �E���Qf����4����L{��8����ȃzY��dx��:��<W�s
(���Gj�M��	�wU�fp��d��EK\L��.��c߶�k���U0�m��t���gx[�t��T�V�&Y�*�5d]����P�5)�1�M:�D�1}5���VpׄE���B�"�+(����Z����ﳩ"w�+<y�q�rf!��\o����m�,���oi��S����.&�)�g�d�y�[9f́�{�&V(�X.�i�Q�m�(���ERZI v�y�S�Y{�n.�%�tg.X�e��y����x�#q8���c��.t2��rJĠ)~�.�x�!ڌ$�AT�!�[v��uז��������5ׇM��F��TA�-���0��ظ�a��%�����hg���6�F�&��Iζ5Zk�<�Ec�������S*�tۮ��x��<.0�upo��y��-ٍ�q�{�!����!��9r]��eڳ���,�8�Y6Q��L�O,�(�&���ګq�xv��<\K3��u�s��KK��x�:���F��/tq��������Z�$E���k��N�NکCs�[��7�8��q�Q�Ǳ�F�e-��������2���B�C�� B��,���u���g���冫]�ה��|�����R��1g.�ڄl��s9�ݏ~q��� v8�ǎ���<D���6�b��j�4�6�VS�#'�]� �;<e�κ�J���g\^�;��7���(��&���I
��iж=/=Ci5��ݷ���=Wj>�\�,�q��w��y��aǙ@���r6�r�UhT�N�M6OR(@i�^9��*�;�L�� �<w�\��4�2@L�3���ڳ�J�<Y��i��ø؋�s�i�����w��R�V� �VVղ�-#��c����lqUj6�{�L4�@���/C��]c��g����.��#s�,g�7�N����W���`�(�Q8�u�l��|�nXGb�w��&�+������%�v��D� �����g5�`�����j�7�Jǋ�`8���]]F��}��-�.�C+��$lPM}%�D�	%�^j���5Oo��G�cn��O3�̳����zO=�s����{�`���*٠��*��垎4|VTd��I*�>�d���ݖ9��zvn����O>���<�hSd�ks��%{4��i��tk��}>�gW�آ!��@Ȩ ໛�PT�S�><y��ѣ�漏�>�zBY��ݫ@w/6(�}�%ER���y}lI6=5ҙ�^�F`>�˹1O��e��dF��)��x��~��Uk�"8�%�����v����\[��ֽ��̈A�|�`PA5��i�����n��V�D�kN�`[-�T�Q���k�V�8c*
*G���Y��k�c�8)k(�>��y�	�ؠ˻��ae!��G�z��6�y ɫ .Ո՘E�\r�,x����c�0��֬�*�Ԣw�UFu�(�]e&H	 &�A��?x�#�-��u$���^=EpN�D���Gm��7&�^����|{͑�����]�m�*�FکW�tۦ޶ȿ"�q�����_����f!��c��$SU�{�G�(�3�ӀK�����Y3�(1��T,���.��t�$��}��r������x��j`·&3� ��A�Q�U�ޑK:����p.#/�A.��^<��Y��ѭ�u��w,�!f�̴�G@���
�*Ě�*͇��Z��^N4��C^Z�Q�$�W��I&nfh�V8	�\t�;k��kB��V��d8w\T����H�,���#6��b��jn]�|qjRgk�6��ψzʭP�9,!d�@�&��\�1-2��ʓ�bR}��fT�e�,wsʯFN�{޳u��r��ϻn��*��'jv �������/�}����[b�rZ�V�e��0�Mi����ϸ<�Wj!6��x�A�0�M�	�����M�P�,������r ͖x�;XI�P<y���;U�(e��	��c"�g3TQe
�n��'��o������m��7u�&�C5 �ZVu�MD4_�x� ���g}3�6�7cT�97j`-�[���� �!mL�����m�}�kĵ�H:�+*r��P���~�Q��e�>� ��Aǹ˩�#1q�֢�&/>��.���[D��-5k.3_n��R����j%5T�Z֚��7�ˡ�������}q\��#��v1rN���/�Ϊ]af��:�ĸn�I�xɸ��ݵ��ғ���Ӝ�Ю��r��6�n����<��M+#yc@��SK�\�q�g�*'tP�x�$n�� �x�/л�q���l�"�I)SS)J����_g�p���㹛��)j�+���:�{���j�O�����xw��g�fec�uj��]؊ǿ!�q�K�e�f��{�-�*�}����*��H������\f�C�ʖL��7G��"���0-�=���;�SѺ�f�oO��=��BY��c�9K2�z��f/��4���-c/��-��[,����K5�TF�Z}�l���J�,���d�i?�E��x�)u�u$6��$Z,c�7*��M��S�r�{��\k|��Z��ߒ��d����TH喒��]ü�{�ޗ�\� ��h:�� w�J���/�����[����h#L]�vS&�Fv�,���K\i92���8�@��2:�@���g�g��{�_$�; ����[�E�aJm���������|}��o��r�0�][ǯڜ5��I�* |�=�g���4D�b���f��t�Aڔ�ieF�e��:n�5��7'%`�Oi�3��>�_MNF�x̘����$� ✪�cS��f&�2�R�MMhS�\�ͪ�l׎Fk/UU �����´ى���9b'��~�������j�J���U\�����Z�]�܆pZ��nZ�ƌϞx�Y���J9E���;�yOi�����	�� �����t�����K������wiPl5�s��7i¢����Y��8�5�о�}ۄ�����9�'����'W�d�cA�E�ն��P�\�I����m8H�LI�p�.wl�!���Q7!�ev�/*�(�F��i˹��6�U�X��!�ظ�Z�j����cx����훧�7~V�'��[�:��BB��`�8�Z����q��<���Oi����p�f����)�7�eo*�¦�<'�e��E��+[�=�G"�r�OO�j��c�Z�v� �|��ш�Ԫ��g'�*���V^����|�*A ����;*�͘s"htĤ@}�����s� q�R����H ggr��_|sejn�?~��4���Ԧ�f�i���xi�����hc{klsg����+����l��k}�}n�]�X���Ȳ������W��X�GD�&u-�E�Y4��)d:���[�Ӻ&f�����$�����ͮ-�F;�����\z��1���;��!Wv��O5�����%��d�g[�P���P�ܣǞ��k�K�i�������Y]��\Q���:)���|^�w��|��U�m.y"�KT��G��fyf��fx 'F��F+l��LSq�X��/�:f�x��{�s��MO5��U�=(�).@��A؇wx����Y؃�����A����ڜ��4�.}�&zP�;�YZ�t�  z�Ț�
�;�1���gWU�<���"���V7�{��� H��,r]�3���XM+�����T�Qpsh�;��*Uxr{��`�>q�3��+i�
��v^4��͇�5�dC���غ� {��Ԋ��}}�� �`)�X&I�h�UkԦ�+�Eۀѳ�[�V�6tݦ��Ȱx����,����4�M�"#�8>�U��=uj�4��+A����ݹ��;)��31ff3E�^��3R�,!�,(hhci���42��8۳�{�:�]��-׎�{б�:�]��C&���Oя���G�\���d��p<� �x��]�i�1@=����Cz�x�XV�T���z9T�G q�Z����ӑ�喻��6@�Y��7Ev�`zivs��N$ <;b�HY�[�fD^m�fe�ɩq�=�e0gZ�~k�6�}�'�qhӒ�H��P$駈�݌9ɖb3$�ڨ���L5�9w�B��'�k��kDNЬ}���s-}]n��
�4ǆc>�6@�3ީn*Tζe�K��I��NJL��4Ī�Fw�x�4�"�۶[�<�|겵���^��܎^����*�;�'�1�*V�N$V��(�����U�� ��Л�@����8vL$��qڠ��u���a=l���X�:�{@��Ǜ��d!����J�4�"��ơ ��g��G�������a�sN�wU�d����`�ȋ9��j>+2�B3���vm���c��Ѷh�\�V,v�v�K`������Zx��e��{TX�;�s����i6#vk���mr`��"�I�Ĕ3><{�q.�e�4�Q����oix�-�WnѴ�ֆ��>�]�y����k���FZu{�>w74iUΰ.�ym���j t��g��d�(� �����3|wY�2�rV���"�N=kbpwϚ�Y=�\�g�dE�5c�t���;�lk#z�x���4�n�n�6ӝ;pB�.rKdLSӅ�`��:���&a�k�`���{%�ٹXq�h�k2��aKS�X4�#	�3L����p�!�J���n�=�N)-
T⟂� OƖ�5�*7���Q��6�z|_a�U�|�Μ����A���9�&�Y����Zd��L�b���t�:���_l�?b$?�K*]9w�2~�p�z�*�G��za��O�U`�r�m"f}�&��	l�p�ϯ^)fUx��O�:���@mcl����ȃ�L\�$ZL�ӱ�>ⵡ�3#)�Nc ��p�QiYw��b��NXl.r��1g�`����{u�-!�g�Д�!���a;�am0�#���>����Q���e5��RZY��e�p�C������ӆ���&�%�� ��E�j���֘�n��rU���5���p��yD8��""������y�<����pԎU���zo(�G��>���܇12�`���S5rj��a�y�T*�������W�4���W���K) N�R1[@	l��l��b}�l���J�@|�libU D��Ǳ�(M+� h�m��^0F�j�p��s��5t�Kc3{��VZ�}�z1|f�X0m+&�*
�����7=�J��ĕ�.]czv�q\)��Jq��I����m'�h��!��lh���Gj��5_��Pn{^�5�w�
eΜ0w�ʷ��,�M.��v1~�i����fǁ�`gn*VȎa�&r��rS)k$R+mz^y���\��~����V`ڛ���M!ݲ�h��cg>����J�}[z�����{Ua��3���ǹF�z���5��t�Y����Z���ej��dP�]�?����>9�3��c�ә�� qr���M��~�� ̴�[�};2�z��U�s���9���:f�q�$v�=���B�$�P���E��[��	If�Z�y�����yK�>x��AǓt�r;S� 6����P��3��ǥ5�tz�dCh@�Qȋ��ڔOV��[�C�Z���w%2EP�0�됒�/4C��4{�^�+�<���9�g���*U�Q޵Ş|�7S�������.�6ck�;kd{T���N�V/�ֶ�UK�-r�+-A���hYf�w3n�CGF�b�0��	�a*�ƫ�b�ѵԙ�Hd�(�[���, a��6m��Smv��_6Ǜ�D��6ƫ�h�&�������*W����Ɓ��&��C��;G��r��,v�H�5��Ğ��w\��f^�Ig�Ѱ�|��,�(ۨ�/��6x|r%������5-�
��0�N���2��g�D����賧(���s
���5�$sg��s�+��"θɁ����F�u6C��3u���p�Za��E�6�ZXU�CÅ�,�v1���p�R�Y�ׁ�;�����f���T,NEb��Nf�֟��'�4�Fm74\x�T_9q�"�s��v� r�8��$Y���M�=��z:�nE���|-um�S@�0U6�1��o(9e� 2\0�Y���B�]�|L�^���S�.~�b�C�=�;����j�U��{^c�uj��?Y����zIF��$��I �� P{�@=��B���߯����L&1@��i����fW�$UE("B""ފT	DEJ��4�@a Q>D r ��"�����
�YgRYq\E(��  cK"�"
a��D���S,�J
Z�b(��[�T�I J��@[E�
��  ��7���B���p
�wE,��;y0��  �(�� �����
�_[L�3�˙�ޅ��7�^������Y�uý����ä���]��Ϭ��74�Ԏ��B矂}=��V������ܟ������A �!���/����S�A �Q懊��o~�>��:���b�B��^{�8����B�������"!8�)^P;?@�pa#�;H3T� *��0�!��d(��i��R�+�<e=OQp���� �/߻��v�sL� �"��@�$B(�"��"��$(�(� �$ ) �E�D�@ 	b�b	b��$@��E AVA`EP�@ ARH�B  DVHXH�`D E�  DVE�@ E0D D@�X�T� D�#�U�U@RRQB1U @T�X @RQ`ERT @�FP�R	dHČ`B�`B`���Q Όy�*���6�l����Ω�Y��@4�0	�#����/`��	� �N�3�j;�E�9����A47����q ���� 9�,<=l�D�p�p�9pg<���f��=�]����.�t>��F<{w���<H�=�� t�H������Ñզ��kކ�s�c�
��b];Q@=���_	�O[h�V�z��	�=F�ä���N!@( ����^���^-,�t����8���2�>%aC�Ɂ�@�˅E� �"�[v�C��О�I�nh� �a=�9� 5��k�5���$I�(�B��>T=���{X�"�QG����4���W�E;�����@9:�?L�f��MS�$0�$`j�_��Y(���l�w��<����x�M.&�w��\�����h����:l^2���A���-OC����4��i� <�ŞM��g�8}f�A�( ������	��&N���u'p�Y��(���������0�s���]�=d@�������&����"�(H��= 